VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_qarma
  CLASS BLOCK ;
  FOREIGN wrapped_qarma ;
  ORIGIN 0.000 0.000 ;
  SIZE 360.000 BY 360.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 356.000 30.270 360.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 1.400 360.000 2.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 95.920 360.000 96.520 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 105.440 360.000 106.040 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 114.960 360.000 115.560 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 123.800 360.000 124.400 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 133.320 360.000 133.920 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 142.840 360.000 143.440 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 152.360 360.000 152.960 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 161.880 360.000 162.480 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 171.400 360.000 172.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 180.920 360.000 181.520 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 10.240 360.000 10.840 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 190.440 360.000 191.040 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 199.960 360.000 200.560 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 209.480 360.000 210.080 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 219.000 360.000 219.600 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 228.520 360.000 229.120 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 238.040 360.000 238.640 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 246.880 360.000 247.480 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 256.400 360.000 257.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 265.920 360.000 266.520 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 275.440 360.000 276.040 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 19.760 360.000 20.360 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 284.960 360.000 285.560 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 294.480 360.000 295.080 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 304.000 360.000 304.600 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 313.520 360.000 314.120 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 323.040 360.000 323.640 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 332.560 360.000 333.160 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 342.080 360.000 342.680 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 351.600 360.000 352.200 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 29.280 360.000 29.880 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 38.800 360.000 39.400 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 48.320 360.000 48.920 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 57.840 360.000 58.440 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 67.360 360.000 67.960 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 76.880 360.000 77.480 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 86.400 360.000 87.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 7.520 360.000 8.120 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 102.040 360.000 102.640 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 111.560 360.000 112.160 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 121.080 360.000 121.680 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 130.600 360.000 131.200 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 140.120 360.000 140.720 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 149.640 360.000 150.240 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 159.160 360.000 159.760 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 168.000 360.000 168.600 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 177.520 360.000 178.120 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 187.040 360.000 187.640 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 17.040 360.000 17.640 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 196.560 360.000 197.160 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 206.080 360.000 206.680 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 215.600 360.000 216.200 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 225.120 360.000 225.720 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 234.640 360.000 235.240 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 244.160 360.000 244.760 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 253.680 360.000 254.280 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 263.200 360.000 263.800 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 272.720 360.000 273.320 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 281.560 360.000 282.160 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 26.560 360.000 27.160 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 291.080 360.000 291.680 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 300.600 360.000 301.200 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 310.120 360.000 310.720 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 319.640 360.000 320.240 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 329.160 360.000 329.760 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 338.680 360.000 339.280 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 348.200 360.000 348.800 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 357.720 360.000 358.320 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 36.080 360.000 36.680 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 44.920 360.000 45.520 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 54.440 360.000 55.040 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 63.960 360.000 64.560 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 73.480 360.000 74.080 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 83.000 360.000 83.600 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 92.520 360.000 93.120 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 4.120 360.000 4.720 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 98.640 360.000 99.240 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 108.160 360.000 108.760 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 117.680 360.000 118.280 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 127.200 360.000 127.800 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 136.720 360.000 137.320 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 146.240 360.000 146.840 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 155.760 360.000 156.360 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 165.280 360.000 165.880 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 174.800 360.000 175.400 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 184.320 360.000 184.920 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 13.640 360.000 14.240 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 193.840 360.000 194.440 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 202.680 360.000 203.280 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 212.200 360.000 212.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 221.720 360.000 222.320 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 231.240 360.000 231.840 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 240.760 360.000 241.360 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 250.280 360.000 250.880 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 259.800 360.000 260.400 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 269.320 360.000 269.920 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 278.840 360.000 279.440 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 23.160 360.000 23.760 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 288.360 360.000 288.960 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 297.880 360.000 298.480 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 307.400 360.000 308.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 316.920 360.000 317.520 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 325.760 360.000 326.360 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 335.280 360.000 335.880 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 344.800 360.000 345.400 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 354.320 360.000 354.920 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 32.680 360.000 33.280 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 42.200 360.000 42.800 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 51.720 360.000 52.320 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 61.240 360.000 61.840 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 70.760 360.000 71.360 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 80.280 360.000 80.880 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 356.000 89.120 360.000 89.720 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 356.000 353.190 360.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 356.000 357.790 360.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 0.000 263.490 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 0.000 202.310 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.720 4.000 239.320 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.160 4.000 244.760 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 283.600 4.000 284.200 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 294.480 4.000 295.080 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.920 4.000 334.520 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END la_oenb[31]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.160 4.000 210.760 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 356.000 34.870 360.000 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 356.000 2.670 360.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 356.000 7.270 360.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 356.000 25.670 360.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 356.000 57.870 360.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 356.000 103.870 360.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 356.000 108.470 360.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 356.000 113.070 360.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 356.000 117.670 360.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 356.000 122.730 360.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 356.000 127.330 360.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 356.000 131.930 360.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 356.000 136.530 360.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 356.000 141.130 360.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 356.000 145.730 360.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 356.000 62.470 360.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 356.000 150.330 360.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 356.000 154.930 360.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 356.000 159.530 360.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 356.000 164.130 360.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 356.000 168.730 360.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 356.000 173.330 360.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 356.000 177.930 360.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 356.000 182.530 360.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 356.000 187.130 360.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 356.000 191.730 360.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 356.000 67.070 360.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 356.000 196.330 360.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 356.000 200.930 360.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 356.000 71.670 360.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 356.000 76.270 360.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 356.000 80.870 360.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 356.000 85.470 360.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 356.000 90.070 360.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 356.000 94.670 360.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 356.000 99.270 360.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 356.000 16.470 360.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 356.000 205.530 360.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 356.000 251.990 360.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 356.000 256.590 360.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 356.000 261.190 360.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 356.000 265.790 360.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 356.000 270.390 360.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 356.000 274.990 360.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 356.000 279.590 360.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 356.000 284.190 360.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 356.000 288.790 360.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 356.000 293.390 360.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 356.000 210.130 360.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 356.000 297.990 360.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 356.000 302.590 360.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 356.000 307.190 360.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 356.000 311.790 360.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 356.000 316.390 360.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 356.000 320.990 360.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 356.000 325.590 360.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 356.000 330.190 360.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 356.000 334.790 360.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 356.000 339.390 360.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 356.000 214.730 360.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 356.000 343.990 360.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 356.000 348.590 360.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 356.000 219.330 360.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 356.000 223.930 360.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 356.000 228.530 360.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 356.000 233.130 360.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 356.000 237.730 360.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 356.000 242.790 360.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 356.000 247.390 360.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 4.000 155.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.280 4.000 165.880 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 356.000 39.470 360.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 356.000 44.070 360.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 356.000 48.670 360.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 356.000 53.270 360.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 356.000 11.870 360.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 356.000 21.070 360.000 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 348.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 348.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 348.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 348.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 348.400 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 348.160 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 348.160 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 348.160 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 348.160 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 348.160 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 348.160 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 348.160 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 348.160 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 348.160 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 348.160 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 348.160 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 348.160 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 348.160 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 348.160 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 348.160 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 354.200 348.245 ;
      LAYER met1 ;
        RECT 2.370 10.640 357.810 352.200 ;
      LAYER met2 ;
        RECT 2.950 355.720 6.710 358.205 ;
        RECT 7.550 355.720 11.310 358.205 ;
        RECT 12.150 355.720 15.910 358.205 ;
        RECT 16.750 355.720 20.510 358.205 ;
        RECT 21.350 355.720 25.110 358.205 ;
        RECT 25.950 355.720 29.710 358.205 ;
        RECT 30.550 355.720 34.310 358.205 ;
        RECT 35.150 355.720 38.910 358.205 ;
        RECT 39.750 355.720 43.510 358.205 ;
        RECT 44.350 355.720 48.110 358.205 ;
        RECT 48.950 355.720 52.710 358.205 ;
        RECT 53.550 355.720 57.310 358.205 ;
        RECT 58.150 355.720 61.910 358.205 ;
        RECT 62.750 355.720 66.510 358.205 ;
        RECT 67.350 355.720 71.110 358.205 ;
        RECT 71.950 355.720 75.710 358.205 ;
        RECT 76.550 355.720 80.310 358.205 ;
        RECT 81.150 355.720 84.910 358.205 ;
        RECT 85.750 355.720 89.510 358.205 ;
        RECT 90.350 355.720 94.110 358.205 ;
        RECT 94.950 355.720 98.710 358.205 ;
        RECT 99.550 355.720 103.310 358.205 ;
        RECT 104.150 355.720 107.910 358.205 ;
        RECT 108.750 355.720 112.510 358.205 ;
        RECT 113.350 355.720 117.110 358.205 ;
        RECT 117.950 355.720 122.170 358.205 ;
        RECT 123.010 355.720 126.770 358.205 ;
        RECT 127.610 355.720 131.370 358.205 ;
        RECT 132.210 355.720 135.970 358.205 ;
        RECT 136.810 355.720 140.570 358.205 ;
        RECT 141.410 355.720 145.170 358.205 ;
        RECT 146.010 355.720 149.770 358.205 ;
        RECT 150.610 355.720 154.370 358.205 ;
        RECT 155.210 355.720 158.970 358.205 ;
        RECT 159.810 355.720 163.570 358.205 ;
        RECT 164.410 355.720 168.170 358.205 ;
        RECT 169.010 355.720 172.770 358.205 ;
        RECT 173.610 355.720 177.370 358.205 ;
        RECT 178.210 355.720 181.970 358.205 ;
        RECT 182.810 355.720 186.570 358.205 ;
        RECT 187.410 355.720 191.170 358.205 ;
        RECT 192.010 355.720 195.770 358.205 ;
        RECT 196.610 355.720 200.370 358.205 ;
        RECT 201.210 355.720 204.970 358.205 ;
        RECT 205.810 355.720 209.570 358.205 ;
        RECT 210.410 355.720 214.170 358.205 ;
        RECT 215.010 355.720 218.770 358.205 ;
        RECT 219.610 355.720 223.370 358.205 ;
        RECT 224.210 355.720 227.970 358.205 ;
        RECT 228.810 355.720 232.570 358.205 ;
        RECT 233.410 355.720 237.170 358.205 ;
        RECT 238.010 355.720 242.230 358.205 ;
        RECT 243.070 355.720 246.830 358.205 ;
        RECT 247.670 355.720 251.430 358.205 ;
        RECT 252.270 355.720 256.030 358.205 ;
        RECT 256.870 355.720 260.630 358.205 ;
        RECT 261.470 355.720 265.230 358.205 ;
        RECT 266.070 355.720 269.830 358.205 ;
        RECT 270.670 355.720 274.430 358.205 ;
        RECT 275.270 355.720 279.030 358.205 ;
        RECT 279.870 355.720 283.630 358.205 ;
        RECT 284.470 355.720 288.230 358.205 ;
        RECT 289.070 355.720 292.830 358.205 ;
        RECT 293.670 355.720 297.430 358.205 ;
        RECT 298.270 355.720 302.030 358.205 ;
        RECT 302.870 355.720 306.630 358.205 ;
        RECT 307.470 355.720 311.230 358.205 ;
        RECT 312.070 355.720 315.830 358.205 ;
        RECT 316.670 355.720 320.430 358.205 ;
        RECT 321.270 355.720 325.030 358.205 ;
        RECT 325.870 355.720 329.630 358.205 ;
        RECT 330.470 355.720 334.230 358.205 ;
        RECT 335.070 355.720 338.830 358.205 ;
        RECT 339.670 355.720 343.430 358.205 ;
        RECT 344.270 355.720 348.030 358.205 ;
        RECT 348.870 355.720 352.630 358.205 ;
        RECT 353.470 355.720 357.230 358.205 ;
        RECT 2.400 4.280 357.780 355.720 ;
        RECT 2.400 1.515 2.570 4.280 ;
        RECT 3.410 1.515 8.090 4.280 ;
        RECT 8.930 1.515 13.610 4.280 ;
        RECT 14.450 1.515 19.130 4.280 ;
        RECT 19.970 1.515 24.650 4.280 ;
        RECT 25.490 1.515 30.170 4.280 ;
        RECT 31.010 1.515 35.690 4.280 ;
        RECT 36.530 1.515 41.210 4.280 ;
        RECT 42.050 1.515 46.730 4.280 ;
        RECT 47.570 1.515 52.250 4.280 ;
        RECT 53.090 1.515 57.770 4.280 ;
        RECT 58.610 1.515 63.290 4.280 ;
        RECT 64.130 1.515 68.810 4.280 ;
        RECT 69.650 1.515 74.330 4.280 ;
        RECT 75.170 1.515 79.850 4.280 ;
        RECT 80.690 1.515 85.370 4.280 ;
        RECT 86.210 1.515 90.890 4.280 ;
        RECT 91.730 1.515 96.410 4.280 ;
        RECT 97.250 1.515 101.930 4.280 ;
        RECT 102.770 1.515 107.450 4.280 ;
        RECT 108.290 1.515 112.970 4.280 ;
        RECT 113.810 1.515 118.490 4.280 ;
        RECT 119.330 1.515 124.470 4.280 ;
        RECT 125.310 1.515 129.990 4.280 ;
        RECT 130.830 1.515 135.510 4.280 ;
        RECT 136.350 1.515 141.030 4.280 ;
        RECT 141.870 1.515 146.550 4.280 ;
        RECT 147.390 1.515 152.070 4.280 ;
        RECT 152.910 1.515 157.590 4.280 ;
        RECT 158.430 1.515 163.110 4.280 ;
        RECT 163.950 1.515 168.630 4.280 ;
        RECT 169.470 1.515 174.150 4.280 ;
        RECT 174.990 1.515 179.670 4.280 ;
        RECT 180.510 1.515 185.190 4.280 ;
        RECT 186.030 1.515 190.710 4.280 ;
        RECT 191.550 1.515 196.230 4.280 ;
        RECT 197.070 1.515 201.750 4.280 ;
        RECT 202.590 1.515 207.270 4.280 ;
        RECT 208.110 1.515 212.790 4.280 ;
        RECT 213.630 1.515 218.310 4.280 ;
        RECT 219.150 1.515 223.830 4.280 ;
        RECT 224.670 1.515 229.350 4.280 ;
        RECT 230.190 1.515 234.870 4.280 ;
        RECT 235.710 1.515 240.390 4.280 ;
        RECT 241.230 1.515 246.370 4.280 ;
        RECT 247.210 1.515 251.890 4.280 ;
        RECT 252.730 1.515 257.410 4.280 ;
        RECT 258.250 1.515 262.930 4.280 ;
        RECT 263.770 1.515 268.450 4.280 ;
        RECT 269.290 1.515 273.970 4.280 ;
        RECT 274.810 1.515 279.490 4.280 ;
        RECT 280.330 1.515 285.010 4.280 ;
        RECT 285.850 1.515 290.530 4.280 ;
        RECT 291.370 1.515 296.050 4.280 ;
        RECT 296.890 1.515 301.570 4.280 ;
        RECT 302.410 1.515 307.090 4.280 ;
        RECT 307.930 1.515 312.610 4.280 ;
        RECT 313.450 1.515 318.130 4.280 ;
        RECT 318.970 1.515 323.650 4.280 ;
        RECT 324.490 1.515 329.170 4.280 ;
        RECT 330.010 1.515 334.690 4.280 ;
        RECT 335.530 1.515 340.210 4.280 ;
        RECT 341.050 1.515 345.730 4.280 ;
        RECT 346.570 1.515 351.250 4.280 ;
        RECT 352.090 1.515 356.770 4.280 ;
        RECT 357.610 1.515 357.780 4.280 ;
      LAYER met3 ;
        RECT 4.000 357.360 355.600 358.185 ;
        RECT 4.400 357.320 355.600 357.360 ;
        RECT 4.400 355.960 356.000 357.320 ;
        RECT 4.000 355.320 356.000 355.960 ;
        RECT 4.000 353.920 355.600 355.320 ;
        RECT 4.000 352.600 356.000 353.920 ;
        RECT 4.000 351.920 355.600 352.600 ;
        RECT 4.400 351.200 355.600 351.920 ;
        RECT 4.400 350.520 356.000 351.200 ;
        RECT 4.000 349.200 356.000 350.520 ;
        RECT 4.000 347.800 355.600 349.200 ;
        RECT 4.000 346.480 356.000 347.800 ;
        RECT 4.400 345.800 356.000 346.480 ;
        RECT 4.400 345.080 355.600 345.800 ;
        RECT 4.000 344.400 355.600 345.080 ;
        RECT 4.000 343.080 356.000 344.400 ;
        RECT 4.000 341.680 355.600 343.080 ;
        RECT 4.000 340.360 356.000 341.680 ;
        RECT 4.400 339.680 356.000 340.360 ;
        RECT 4.400 338.960 355.600 339.680 ;
        RECT 4.000 338.280 355.600 338.960 ;
        RECT 4.000 336.280 356.000 338.280 ;
        RECT 4.000 334.920 355.600 336.280 ;
        RECT 4.400 334.880 355.600 334.920 ;
        RECT 4.400 333.560 356.000 334.880 ;
        RECT 4.400 333.520 355.600 333.560 ;
        RECT 4.000 332.160 355.600 333.520 ;
        RECT 4.000 330.160 356.000 332.160 ;
        RECT 4.000 329.480 355.600 330.160 ;
        RECT 4.400 328.760 355.600 329.480 ;
        RECT 4.400 328.080 356.000 328.760 ;
        RECT 4.000 326.760 356.000 328.080 ;
        RECT 4.000 325.360 355.600 326.760 ;
        RECT 4.000 324.040 356.000 325.360 ;
        RECT 4.400 322.640 355.600 324.040 ;
        RECT 4.000 320.640 356.000 322.640 ;
        RECT 4.000 319.240 355.600 320.640 ;
        RECT 4.000 317.920 356.000 319.240 ;
        RECT 4.400 316.520 355.600 317.920 ;
        RECT 4.000 314.520 356.000 316.520 ;
        RECT 4.000 313.120 355.600 314.520 ;
        RECT 4.000 312.480 356.000 313.120 ;
        RECT 4.400 311.120 356.000 312.480 ;
        RECT 4.400 311.080 355.600 311.120 ;
        RECT 4.000 309.720 355.600 311.080 ;
        RECT 4.000 308.400 356.000 309.720 ;
        RECT 4.000 307.040 355.600 308.400 ;
        RECT 4.400 307.000 355.600 307.040 ;
        RECT 4.400 305.640 356.000 307.000 ;
        RECT 4.000 305.000 356.000 305.640 ;
        RECT 4.000 303.600 355.600 305.000 ;
        RECT 4.000 301.600 356.000 303.600 ;
        RECT 4.400 300.200 355.600 301.600 ;
        RECT 4.000 298.880 356.000 300.200 ;
        RECT 4.000 297.480 355.600 298.880 ;
        RECT 4.000 295.480 356.000 297.480 ;
        RECT 4.400 294.080 355.600 295.480 ;
        RECT 4.000 292.080 356.000 294.080 ;
        RECT 4.000 290.680 355.600 292.080 ;
        RECT 4.000 290.040 356.000 290.680 ;
        RECT 4.400 289.360 356.000 290.040 ;
        RECT 4.400 288.640 355.600 289.360 ;
        RECT 4.000 287.960 355.600 288.640 ;
        RECT 4.000 285.960 356.000 287.960 ;
        RECT 4.000 284.600 355.600 285.960 ;
        RECT 4.400 284.560 355.600 284.600 ;
        RECT 4.400 283.200 356.000 284.560 ;
        RECT 4.000 282.560 356.000 283.200 ;
        RECT 4.000 281.160 355.600 282.560 ;
        RECT 4.000 279.840 356.000 281.160 ;
        RECT 4.000 279.160 355.600 279.840 ;
        RECT 4.400 278.440 355.600 279.160 ;
        RECT 4.400 277.760 356.000 278.440 ;
        RECT 4.000 276.440 356.000 277.760 ;
        RECT 4.000 275.040 355.600 276.440 ;
        RECT 4.000 273.720 356.000 275.040 ;
        RECT 4.000 273.040 355.600 273.720 ;
        RECT 4.400 272.320 355.600 273.040 ;
        RECT 4.400 271.640 356.000 272.320 ;
        RECT 4.000 270.320 356.000 271.640 ;
        RECT 4.000 268.920 355.600 270.320 ;
        RECT 4.000 267.600 356.000 268.920 ;
        RECT 4.400 266.920 356.000 267.600 ;
        RECT 4.400 266.200 355.600 266.920 ;
        RECT 4.000 265.520 355.600 266.200 ;
        RECT 4.000 264.200 356.000 265.520 ;
        RECT 4.000 262.800 355.600 264.200 ;
        RECT 4.000 262.160 356.000 262.800 ;
        RECT 4.400 260.800 356.000 262.160 ;
        RECT 4.400 260.760 355.600 260.800 ;
        RECT 4.000 259.400 355.600 260.760 ;
        RECT 4.000 257.400 356.000 259.400 ;
        RECT 4.000 256.040 355.600 257.400 ;
        RECT 4.400 256.000 355.600 256.040 ;
        RECT 4.400 254.680 356.000 256.000 ;
        RECT 4.400 254.640 355.600 254.680 ;
        RECT 4.000 253.280 355.600 254.640 ;
        RECT 4.000 251.280 356.000 253.280 ;
        RECT 4.000 250.600 355.600 251.280 ;
        RECT 4.400 249.880 355.600 250.600 ;
        RECT 4.400 249.200 356.000 249.880 ;
        RECT 4.000 247.880 356.000 249.200 ;
        RECT 4.000 246.480 355.600 247.880 ;
        RECT 4.000 245.160 356.000 246.480 ;
        RECT 4.400 243.760 355.600 245.160 ;
        RECT 4.000 241.760 356.000 243.760 ;
        RECT 4.000 240.360 355.600 241.760 ;
        RECT 4.000 239.720 356.000 240.360 ;
        RECT 4.400 239.040 356.000 239.720 ;
        RECT 4.400 238.320 355.600 239.040 ;
        RECT 4.000 237.640 355.600 238.320 ;
        RECT 4.000 235.640 356.000 237.640 ;
        RECT 4.000 234.240 355.600 235.640 ;
        RECT 4.000 233.600 356.000 234.240 ;
        RECT 4.400 232.240 356.000 233.600 ;
        RECT 4.400 232.200 355.600 232.240 ;
        RECT 4.000 230.840 355.600 232.200 ;
        RECT 4.000 229.520 356.000 230.840 ;
        RECT 4.000 228.160 355.600 229.520 ;
        RECT 4.400 228.120 355.600 228.160 ;
        RECT 4.400 226.760 356.000 228.120 ;
        RECT 4.000 226.120 356.000 226.760 ;
        RECT 4.000 224.720 355.600 226.120 ;
        RECT 4.000 222.720 356.000 224.720 ;
        RECT 4.400 221.320 355.600 222.720 ;
        RECT 4.000 220.000 356.000 221.320 ;
        RECT 4.000 218.600 355.600 220.000 ;
        RECT 4.000 217.280 356.000 218.600 ;
        RECT 4.400 216.600 356.000 217.280 ;
        RECT 4.400 215.880 355.600 216.600 ;
        RECT 4.000 215.200 355.600 215.880 ;
        RECT 4.000 213.200 356.000 215.200 ;
        RECT 4.000 211.800 355.600 213.200 ;
        RECT 4.000 211.160 356.000 211.800 ;
        RECT 4.400 210.480 356.000 211.160 ;
        RECT 4.400 209.760 355.600 210.480 ;
        RECT 4.000 209.080 355.600 209.760 ;
        RECT 4.000 207.080 356.000 209.080 ;
        RECT 4.000 205.720 355.600 207.080 ;
        RECT 4.400 205.680 355.600 205.720 ;
        RECT 4.400 204.320 356.000 205.680 ;
        RECT 4.000 203.680 356.000 204.320 ;
        RECT 4.000 202.280 355.600 203.680 ;
        RECT 4.000 200.960 356.000 202.280 ;
        RECT 4.000 200.280 355.600 200.960 ;
        RECT 4.400 199.560 355.600 200.280 ;
        RECT 4.400 198.880 356.000 199.560 ;
        RECT 4.000 197.560 356.000 198.880 ;
        RECT 4.000 196.160 355.600 197.560 ;
        RECT 4.000 194.840 356.000 196.160 ;
        RECT 4.400 193.440 355.600 194.840 ;
        RECT 4.000 191.440 356.000 193.440 ;
        RECT 4.000 190.040 355.600 191.440 ;
        RECT 4.000 188.720 356.000 190.040 ;
        RECT 4.400 188.040 356.000 188.720 ;
        RECT 4.400 187.320 355.600 188.040 ;
        RECT 4.000 186.640 355.600 187.320 ;
        RECT 4.000 185.320 356.000 186.640 ;
        RECT 4.000 183.920 355.600 185.320 ;
        RECT 4.000 183.280 356.000 183.920 ;
        RECT 4.400 181.920 356.000 183.280 ;
        RECT 4.400 181.880 355.600 181.920 ;
        RECT 4.000 180.520 355.600 181.880 ;
        RECT 4.000 178.520 356.000 180.520 ;
        RECT 4.000 177.840 355.600 178.520 ;
        RECT 4.400 177.120 355.600 177.840 ;
        RECT 4.400 176.440 356.000 177.120 ;
        RECT 4.000 175.800 356.000 176.440 ;
        RECT 4.000 174.400 355.600 175.800 ;
        RECT 4.000 172.400 356.000 174.400 ;
        RECT 4.000 171.720 355.600 172.400 ;
        RECT 4.400 171.000 355.600 171.720 ;
        RECT 4.400 170.320 356.000 171.000 ;
        RECT 4.000 169.000 356.000 170.320 ;
        RECT 4.000 167.600 355.600 169.000 ;
        RECT 4.000 166.280 356.000 167.600 ;
        RECT 4.400 164.880 355.600 166.280 ;
        RECT 4.000 162.880 356.000 164.880 ;
        RECT 4.000 161.480 355.600 162.880 ;
        RECT 4.000 160.840 356.000 161.480 ;
        RECT 4.400 160.160 356.000 160.840 ;
        RECT 4.400 159.440 355.600 160.160 ;
        RECT 4.000 158.760 355.600 159.440 ;
        RECT 4.000 156.760 356.000 158.760 ;
        RECT 4.000 155.400 355.600 156.760 ;
        RECT 4.400 155.360 355.600 155.400 ;
        RECT 4.400 154.000 356.000 155.360 ;
        RECT 4.000 153.360 356.000 154.000 ;
        RECT 4.000 151.960 355.600 153.360 ;
        RECT 4.000 150.640 356.000 151.960 ;
        RECT 4.000 149.280 355.600 150.640 ;
        RECT 4.400 149.240 355.600 149.280 ;
        RECT 4.400 147.880 356.000 149.240 ;
        RECT 4.000 147.240 356.000 147.880 ;
        RECT 4.000 145.840 355.600 147.240 ;
        RECT 4.000 143.840 356.000 145.840 ;
        RECT 4.400 142.440 355.600 143.840 ;
        RECT 4.000 141.120 356.000 142.440 ;
        RECT 4.000 139.720 355.600 141.120 ;
        RECT 4.000 138.400 356.000 139.720 ;
        RECT 4.400 137.720 356.000 138.400 ;
        RECT 4.400 137.000 355.600 137.720 ;
        RECT 4.000 136.320 355.600 137.000 ;
        RECT 4.000 134.320 356.000 136.320 ;
        RECT 4.000 132.960 355.600 134.320 ;
        RECT 4.400 132.920 355.600 132.960 ;
        RECT 4.400 131.600 356.000 132.920 ;
        RECT 4.400 131.560 355.600 131.600 ;
        RECT 4.000 130.200 355.600 131.560 ;
        RECT 4.000 128.200 356.000 130.200 ;
        RECT 4.000 126.840 355.600 128.200 ;
        RECT 4.400 126.800 355.600 126.840 ;
        RECT 4.400 125.440 356.000 126.800 ;
        RECT 4.000 124.800 356.000 125.440 ;
        RECT 4.000 123.400 355.600 124.800 ;
        RECT 4.000 122.080 356.000 123.400 ;
        RECT 4.000 121.400 355.600 122.080 ;
        RECT 4.400 120.680 355.600 121.400 ;
        RECT 4.400 120.000 356.000 120.680 ;
        RECT 4.000 118.680 356.000 120.000 ;
        RECT 4.000 117.280 355.600 118.680 ;
        RECT 4.000 115.960 356.000 117.280 ;
        RECT 4.400 114.560 355.600 115.960 ;
        RECT 4.000 112.560 356.000 114.560 ;
        RECT 4.000 111.160 355.600 112.560 ;
        RECT 4.000 110.520 356.000 111.160 ;
        RECT 4.400 109.160 356.000 110.520 ;
        RECT 4.400 109.120 355.600 109.160 ;
        RECT 4.000 107.760 355.600 109.120 ;
        RECT 4.000 106.440 356.000 107.760 ;
        RECT 4.000 105.040 355.600 106.440 ;
        RECT 4.000 104.400 356.000 105.040 ;
        RECT 4.400 103.040 356.000 104.400 ;
        RECT 4.400 103.000 355.600 103.040 ;
        RECT 4.000 101.640 355.600 103.000 ;
        RECT 4.000 99.640 356.000 101.640 ;
        RECT 4.000 98.960 355.600 99.640 ;
        RECT 4.400 98.240 355.600 98.960 ;
        RECT 4.400 97.560 356.000 98.240 ;
        RECT 4.000 96.920 356.000 97.560 ;
        RECT 4.000 95.520 355.600 96.920 ;
        RECT 4.000 93.520 356.000 95.520 ;
        RECT 4.400 92.120 355.600 93.520 ;
        RECT 4.000 90.120 356.000 92.120 ;
        RECT 4.000 88.720 355.600 90.120 ;
        RECT 4.000 87.400 356.000 88.720 ;
        RECT 4.400 86.000 355.600 87.400 ;
        RECT 4.000 84.000 356.000 86.000 ;
        RECT 4.000 82.600 355.600 84.000 ;
        RECT 4.000 81.960 356.000 82.600 ;
        RECT 4.400 81.280 356.000 81.960 ;
        RECT 4.400 80.560 355.600 81.280 ;
        RECT 4.000 79.880 355.600 80.560 ;
        RECT 4.000 77.880 356.000 79.880 ;
        RECT 4.000 76.520 355.600 77.880 ;
        RECT 4.400 76.480 355.600 76.520 ;
        RECT 4.400 75.120 356.000 76.480 ;
        RECT 4.000 74.480 356.000 75.120 ;
        RECT 4.000 73.080 355.600 74.480 ;
        RECT 4.000 71.760 356.000 73.080 ;
        RECT 4.000 71.080 355.600 71.760 ;
        RECT 4.400 70.360 355.600 71.080 ;
        RECT 4.400 69.680 356.000 70.360 ;
        RECT 4.000 68.360 356.000 69.680 ;
        RECT 4.000 66.960 355.600 68.360 ;
        RECT 4.000 64.960 356.000 66.960 ;
        RECT 4.400 63.560 355.600 64.960 ;
        RECT 4.000 62.240 356.000 63.560 ;
        RECT 4.000 60.840 355.600 62.240 ;
        RECT 4.000 59.520 356.000 60.840 ;
        RECT 4.400 58.840 356.000 59.520 ;
        RECT 4.400 58.120 355.600 58.840 ;
        RECT 4.000 57.440 355.600 58.120 ;
        RECT 4.000 55.440 356.000 57.440 ;
        RECT 4.000 54.080 355.600 55.440 ;
        RECT 4.400 54.040 355.600 54.080 ;
        RECT 4.400 52.720 356.000 54.040 ;
        RECT 4.400 52.680 355.600 52.720 ;
        RECT 4.000 51.320 355.600 52.680 ;
        RECT 4.000 49.320 356.000 51.320 ;
        RECT 4.000 48.640 355.600 49.320 ;
        RECT 4.400 47.920 355.600 48.640 ;
        RECT 4.400 47.240 356.000 47.920 ;
        RECT 4.000 45.920 356.000 47.240 ;
        RECT 4.000 44.520 355.600 45.920 ;
        RECT 4.000 43.200 356.000 44.520 ;
        RECT 4.000 42.520 355.600 43.200 ;
        RECT 4.400 41.800 355.600 42.520 ;
        RECT 4.400 41.120 356.000 41.800 ;
        RECT 4.000 39.800 356.000 41.120 ;
        RECT 4.000 38.400 355.600 39.800 ;
        RECT 4.000 37.080 356.000 38.400 ;
        RECT 4.400 35.680 355.600 37.080 ;
        RECT 4.000 33.680 356.000 35.680 ;
        RECT 4.000 32.280 355.600 33.680 ;
        RECT 4.000 31.640 356.000 32.280 ;
        RECT 4.400 30.280 356.000 31.640 ;
        RECT 4.400 30.240 355.600 30.280 ;
        RECT 4.000 28.880 355.600 30.240 ;
        RECT 4.000 27.560 356.000 28.880 ;
        RECT 4.000 26.200 355.600 27.560 ;
        RECT 4.400 26.160 355.600 26.200 ;
        RECT 4.400 24.800 356.000 26.160 ;
        RECT 4.000 24.160 356.000 24.800 ;
        RECT 4.000 22.760 355.600 24.160 ;
        RECT 4.000 20.760 356.000 22.760 ;
        RECT 4.000 20.080 355.600 20.760 ;
        RECT 4.400 19.360 355.600 20.080 ;
        RECT 4.400 18.680 356.000 19.360 ;
        RECT 4.000 18.040 356.000 18.680 ;
        RECT 4.000 16.640 355.600 18.040 ;
        RECT 4.000 14.640 356.000 16.640 ;
        RECT 4.400 13.240 355.600 14.640 ;
        RECT 4.000 11.240 356.000 13.240 ;
        RECT 4.000 9.840 355.600 11.240 ;
        RECT 4.000 9.200 356.000 9.840 ;
        RECT 4.400 8.520 356.000 9.200 ;
        RECT 4.400 7.800 355.600 8.520 ;
        RECT 4.000 7.120 355.600 7.800 ;
        RECT 4.000 5.120 356.000 7.120 ;
        RECT 4.000 3.760 355.600 5.120 ;
        RECT 4.400 3.720 355.600 3.760 ;
        RECT 4.400 2.400 356.000 3.720 ;
        RECT 4.400 2.360 355.600 2.400 ;
        RECT 4.000 1.535 355.600 2.360 ;
      LAYER met4 ;
        RECT 26.975 50.495 27.240 328.265 ;
        RECT 29.640 50.495 30.540 328.265 ;
        RECT 32.940 50.495 97.440 328.265 ;
        RECT 99.840 50.495 100.740 328.265 ;
        RECT 103.140 50.495 104.040 328.265 ;
        RECT 106.440 50.495 107.340 328.265 ;
        RECT 109.740 50.495 174.240 328.265 ;
        RECT 176.640 50.495 177.540 328.265 ;
        RECT 179.940 50.495 180.840 328.265 ;
        RECT 183.240 50.495 184.140 328.265 ;
        RECT 186.540 50.495 251.040 328.265 ;
        RECT 253.440 50.495 254.340 328.265 ;
        RECT 256.740 50.495 257.640 328.265 ;
        RECT 260.040 50.495 260.940 328.265 ;
        RECT 263.340 50.495 327.840 328.265 ;
        RECT 330.240 50.495 330.905 328.265 ;
  END
END wrapped_qarma
END LIBRARY

