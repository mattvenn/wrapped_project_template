VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_quad_pwm_fet_drivers
  CLASS BLOCK ;
  FOREIGN wrapped_quad_pwm_fet_drivers ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.790 296.000 25.350 300.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 0.420 300.000 1.620 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 78.620 300.000 79.820 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 86.100 300.000 87.300 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 94.260 300.000 95.460 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 101.740 300.000 102.940 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 109.900 300.000 111.100 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 117.380 300.000 118.580 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 125.540 300.000 126.740 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 133.020 300.000 134.220 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 141.180 300.000 142.380 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 148.660 300.000 149.860 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 7.900 300.000 9.100 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 156.820 300.000 158.020 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 164.300 300.000 165.500 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 172.460 300.000 173.660 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 179.940 300.000 181.140 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 188.100 300.000 189.300 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 195.580 300.000 196.780 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 203.740 300.000 204.940 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 211.220 300.000 212.420 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 219.380 300.000 220.580 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 226.860 300.000 228.060 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 16.060 300.000 17.260 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 235.020 300.000 236.220 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 242.500 300.000 243.700 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 250.660 300.000 251.860 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 258.140 300.000 259.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 266.300 300.000 267.500 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 273.780 300.000 274.980 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 281.940 300.000 283.140 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 289.420 300.000 290.620 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 23.540 300.000 24.740 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 31.700 300.000 32.900 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 39.180 300.000 40.380 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 47.340 300.000 48.540 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 54.820 300.000 56.020 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 62.980 300.000 64.180 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 70.460 300.000 71.660 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 5.180 300.000 6.380 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 83.380 300.000 84.580 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 91.540 300.000 92.740 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 99.020 300.000 100.220 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 107.180 300.000 108.380 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 114.660 300.000 115.860 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 122.820 300.000 124.020 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 130.300 300.000 131.500 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 138.460 300.000 139.660 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 145.940 300.000 147.140 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 154.100 300.000 155.300 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 13.340 300.000 14.540 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 161.580 300.000 162.780 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 169.740 300.000 170.940 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 177.220 300.000 178.420 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 185.380 300.000 186.580 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 192.860 300.000 194.060 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 201.020 300.000 202.220 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 208.500 300.000 209.700 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 216.660 300.000 217.860 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 224.140 300.000 225.340 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 232.300 300.000 233.500 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 20.820 300.000 22.020 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 239.780 300.000 240.980 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 247.940 300.000 249.140 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 255.420 300.000 256.620 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 263.580 300.000 264.780 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 271.060 300.000 272.260 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 279.220 300.000 280.420 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 286.700 300.000 287.900 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 294.860 300.000 296.060 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 28.980 300.000 30.180 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 36.460 300.000 37.660 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 44.620 300.000 45.820 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 52.100 300.000 53.300 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 60.260 300.000 61.460 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 67.740 300.000 68.940 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 75.900 300.000 77.100 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 2.460 300.000 3.660 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 80.660 300.000 81.860 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 88.820 300.000 90.020 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 96.300 300.000 97.500 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 104.460 300.000 105.660 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 111.940 300.000 113.140 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 120.100 300.000 121.300 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 127.580 300.000 128.780 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 135.740 300.000 136.940 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 143.220 300.000 144.420 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 151.380 300.000 152.580 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 10.620 300.000 11.820 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 158.860 300.000 160.060 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 167.020 300.000 168.220 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 174.500 300.000 175.700 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 182.660 300.000 183.860 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 190.140 300.000 191.340 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 198.300 300.000 199.500 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 205.780 300.000 206.980 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 213.940 300.000 215.140 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 221.420 300.000 222.620 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 229.580 300.000 230.780 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 18.100 300.000 19.300 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 237.060 300.000 238.260 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 245.220 300.000 246.420 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 252.700 300.000 253.900 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 260.860 300.000 262.060 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 268.340 300.000 269.540 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 276.500 300.000 277.700 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 283.980 300.000 285.180 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 292.140 300.000 293.340 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 26.260 300.000 27.460 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 33.740 300.000 34.940 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 41.900 300.000 43.100 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 49.380 300.000 50.580 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 57.540 300.000 58.740 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 65.020 300.000 66.220 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 73.180 300.000 74.380 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 297.580 300.000 298.780 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.110 0.000 297.670 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.570 296.000 298.130 300.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.250 0.000 2.810 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.250 0.000 48.810 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.850 0.000 53.410 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.450 0.000 58.010 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.050 0.000 62.610 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.650 0.000 67.210 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.250 0.000 71.810 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.850 0.000 76.410 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.450 0.000 81.010 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.050 0.000 85.610 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.650 0.000 90.210 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.850 0.000 7.410 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.250 0.000 94.810 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.850 0.000 99.410 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.450 0.000 104.010 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.050 0.000 108.610 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.650 0.000 113.210 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.250 0.000 117.810 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.850 0.000 122.410 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450 0.000 127.010 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.050 0.000 131.610 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.650 0.000 136.210 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.450 0.000 12.010 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.250 0.000 140.810 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.850 0.000 145.410 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.050 0.000 16.610 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.650 0.000 21.210 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.250 0.000 25.810 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.850 0.000 30.410 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.450 0.000 35.010 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.050 0.000 39.610 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 0.000 44.210 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.450 0.000 150.010 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.910 0.000 196.470 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.510 0.000 201.070 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.110 0.000 205.670 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.710 0.000 210.270 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.310 0.000 214.870 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.910 0.000 219.470 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.510 0.000 224.070 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.110 0.000 228.670 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.710 0.000 233.270 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.310 0.000 237.870 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.510 0.000 155.070 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.910 0.000 242.470 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.510 0.000 247.070 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.110 0.000 251.670 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.710 0.000 256.270 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.310 0.000 260.870 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.910 0.000 265.470 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.510 0.000 270.070 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.110 0.000 274.670 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.710 0.000 279.270 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.310 0.000 283.870 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.110 0.000 159.670 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.910 0.000 288.470 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.510 0.000 293.070 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.710 0.000 164.270 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.310 0.000 168.870 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.910 0.000 173.470 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.510 0.000 178.070 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.110 0.000 182.670 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.710 0.000 187.270 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.310 0.000 191.870 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.380 4.000 152.580 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.300 4.000 199.500 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.060 4.000 204.260 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.820 4.000 209.020 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.580 4.000 213.780 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.660 4.000 217.860 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.420 4.000 222.620 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.180 4.000 227.380 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.940 4.000 232.140 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.700 4.000 236.900 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.460 4.000 241.660 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.140 4.000 157.340 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.220 4.000 246.420 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.980 4.000 251.180 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.740 4.000 255.940 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.820 4.000 260.020 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.580 4.000 264.780 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.340 4.000 269.540 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.100 4.000 274.300 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.860 4.000 279.060 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.620 4.000 283.820 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.380 4.000 288.580 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.900 4.000 162.100 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.140 4.000 293.340 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.900 4.000 298.100 ;
    END
  END la_oenb[31]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.660 4.000 166.860 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.420 4.000 171.620 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.500 4.000 175.700 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.260 4.000 180.460 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.020 4.000 185.220 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.780 4.000 189.980 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.540 4.000 194.740 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.930 296.000 29.490 300.000 ;
    END
  END user_clock2
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.790 296.000 2.350 300.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.470 296.000 6.030 300.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.110 296.000 21.670 300.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.250 296.000 48.810 300.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.350 296.000 87.910 300.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 296.000 91.590 300.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.170 296.000 95.730 300.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.850 296.000 99.410 300.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 296.000 103.550 300.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.670 296.000 107.230 300.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.810 296.000 111.370 300.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.490 296.000 115.050 300.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.630 296.000 119.190 300.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.310 296.000 122.870 300.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.390 296.000 52.950 300.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.990 296.000 126.550 300.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.130 296.000 130.690 300.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.810 296.000 134.370 300.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.950 296.000 138.510 300.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.630 296.000 142.190 300.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.770 296.000 146.330 300.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.450 296.000 150.010 300.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.590 296.000 154.150 300.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.270 296.000 157.830 300.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.410 296.000 161.970 300.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.070 296.000 56.630 300.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.090 296.000 165.650 300.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.230 296.000 169.790 300.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.210 296.000 60.770 300.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.890 296.000 64.450 300.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 296.000 68.130 300.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.710 296.000 72.270 300.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.390 296.000 75.950 300.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.530 296.000 80.090 300.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.210 296.000 83.770 300.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.290 296.000 13.850 300.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.910 296.000 173.470 300.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.010 296.000 212.570 300.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.690 296.000 216.250 300.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.830 296.000 220.390 300.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.510 296.000 224.070 300.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.650 296.000 228.210 300.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.330 296.000 231.890 300.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.470 296.000 236.030 300.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.150 296.000 239.710 300.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.830 296.000 243.390 300.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.970 296.000 247.530 300.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.050 296.000 177.610 300.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.650 296.000 251.210 300.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.790 296.000 255.350 300.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.470 296.000 259.030 300.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.610 296.000 263.170 300.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.290 296.000 266.850 300.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.430 296.000 270.990 300.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.110 296.000 274.670 300.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.250 296.000 278.810 300.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.930 296.000 282.490 300.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.070 296.000 286.630 300.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.730 296.000 181.290 300.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.750 296.000 290.310 300.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.890 296.000 294.450 300.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.410 296.000 184.970 300.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.550 296.000 189.110 300.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.230 296.000 192.790 300.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.370 296.000 196.930 300.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.050 296.000 200.610 300.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.190 296.000 204.750 300.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.870 296.000 208.430 300.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.780 4.000 2.980 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.020 4.000 49.220 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.780 4.000 53.980 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.540 4.000 58.740 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.300 4.000 63.500 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.060 4.000 68.260 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.820 4.000 73.020 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.580 4.000 77.780 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.340 4.000 82.540 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.100 4.000 87.300 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.180 4.000 91.380 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.860 4.000 7.060 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.940 4.000 96.140 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.700 4.000 100.900 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.460 4.000 105.660 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.220 4.000 110.420 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.980 4.000 115.180 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.740 4.000 119.940 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.500 4.000 124.700 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.260 4.000 129.460 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.340 4.000 133.540 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.100 4.000 138.300 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.620 4.000 11.820 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.860 4.000 143.060 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.620 4.000 147.820 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.380 4.000 16.580 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.140 4.000 21.340 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.900 4.000 26.100 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.660 4.000 30.860 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.420 4.000 35.620 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.180 4.000 40.380 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.940 4.000 45.140 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.610 296.000 33.170 300.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.750 296.000 37.310 300.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 296.000 40.990 300.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.570 296.000 45.130 300.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.150 296.000 9.710 300.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.970 296.000 17.530 300.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 295.635 288.405 ;
      LAYER met1 ;
        RECT 1.910 6.160 298.010 288.560 ;
      LAYER met2 ;
        RECT 2.630 295.720 5.190 298.365 ;
        RECT 6.310 295.720 8.870 298.365 ;
        RECT 9.990 295.720 13.010 298.365 ;
        RECT 14.130 295.720 16.690 298.365 ;
        RECT 17.810 295.720 20.830 298.365 ;
        RECT 21.950 295.720 24.510 298.365 ;
        RECT 25.630 295.720 28.650 298.365 ;
        RECT 29.770 295.720 32.330 298.365 ;
        RECT 33.450 295.720 36.470 298.365 ;
        RECT 37.590 295.720 40.150 298.365 ;
        RECT 41.270 295.720 44.290 298.365 ;
        RECT 45.410 295.720 47.970 298.365 ;
        RECT 49.090 295.720 52.110 298.365 ;
        RECT 53.230 295.720 55.790 298.365 ;
        RECT 56.910 295.720 59.930 298.365 ;
        RECT 61.050 295.720 63.610 298.365 ;
        RECT 64.730 295.720 67.290 298.365 ;
        RECT 68.410 295.720 71.430 298.365 ;
        RECT 72.550 295.720 75.110 298.365 ;
        RECT 76.230 295.720 79.250 298.365 ;
        RECT 80.370 295.720 82.930 298.365 ;
        RECT 84.050 295.720 87.070 298.365 ;
        RECT 88.190 295.720 90.750 298.365 ;
        RECT 91.870 295.720 94.890 298.365 ;
        RECT 96.010 295.720 98.570 298.365 ;
        RECT 99.690 295.720 102.710 298.365 ;
        RECT 103.830 295.720 106.390 298.365 ;
        RECT 107.510 295.720 110.530 298.365 ;
        RECT 111.650 295.720 114.210 298.365 ;
        RECT 115.330 295.720 118.350 298.365 ;
        RECT 119.470 295.720 122.030 298.365 ;
        RECT 123.150 295.720 125.710 298.365 ;
        RECT 126.830 295.720 129.850 298.365 ;
        RECT 130.970 295.720 133.530 298.365 ;
        RECT 134.650 295.720 137.670 298.365 ;
        RECT 138.790 295.720 141.350 298.365 ;
        RECT 142.470 295.720 145.490 298.365 ;
        RECT 146.610 295.720 149.170 298.365 ;
        RECT 150.290 295.720 153.310 298.365 ;
        RECT 154.430 295.720 156.990 298.365 ;
        RECT 158.110 295.720 161.130 298.365 ;
        RECT 162.250 295.720 164.810 298.365 ;
        RECT 165.930 295.720 168.950 298.365 ;
        RECT 170.070 295.720 172.630 298.365 ;
        RECT 173.750 295.720 176.770 298.365 ;
        RECT 177.890 295.720 180.450 298.365 ;
        RECT 181.570 295.720 184.130 298.365 ;
        RECT 185.250 295.720 188.270 298.365 ;
        RECT 189.390 295.720 191.950 298.365 ;
        RECT 193.070 295.720 196.090 298.365 ;
        RECT 197.210 295.720 199.770 298.365 ;
        RECT 200.890 295.720 203.910 298.365 ;
        RECT 205.030 295.720 207.590 298.365 ;
        RECT 208.710 295.720 211.730 298.365 ;
        RECT 212.850 295.720 215.410 298.365 ;
        RECT 216.530 295.720 219.550 298.365 ;
        RECT 220.670 295.720 223.230 298.365 ;
        RECT 224.350 295.720 227.370 298.365 ;
        RECT 228.490 295.720 231.050 298.365 ;
        RECT 232.170 295.720 235.190 298.365 ;
        RECT 236.310 295.720 238.870 298.365 ;
        RECT 239.990 295.720 242.550 298.365 ;
        RECT 243.670 295.720 246.690 298.365 ;
        RECT 247.810 295.720 250.370 298.365 ;
        RECT 251.490 295.720 254.510 298.365 ;
        RECT 255.630 295.720 258.190 298.365 ;
        RECT 259.310 295.720 262.330 298.365 ;
        RECT 263.450 295.720 266.010 298.365 ;
        RECT 267.130 295.720 270.150 298.365 ;
        RECT 271.270 295.720 273.830 298.365 ;
        RECT 274.950 295.720 277.970 298.365 ;
        RECT 279.090 295.720 281.650 298.365 ;
        RECT 282.770 295.720 285.790 298.365 ;
        RECT 286.910 295.720 289.470 298.365 ;
        RECT 290.590 295.720 293.610 298.365 ;
        RECT 294.730 295.720 297.290 298.365 ;
        RECT 1.940 4.280 297.980 295.720 ;
        RECT 1.940 2.195 1.970 4.280 ;
        RECT 3.090 2.195 6.570 4.280 ;
        RECT 7.690 2.195 11.170 4.280 ;
        RECT 12.290 2.195 15.770 4.280 ;
        RECT 16.890 2.195 20.370 4.280 ;
        RECT 21.490 2.195 24.970 4.280 ;
        RECT 26.090 2.195 29.570 4.280 ;
        RECT 30.690 2.195 34.170 4.280 ;
        RECT 35.290 2.195 38.770 4.280 ;
        RECT 39.890 2.195 43.370 4.280 ;
        RECT 44.490 2.195 47.970 4.280 ;
        RECT 49.090 2.195 52.570 4.280 ;
        RECT 53.690 2.195 57.170 4.280 ;
        RECT 58.290 2.195 61.770 4.280 ;
        RECT 62.890 2.195 66.370 4.280 ;
        RECT 67.490 2.195 70.970 4.280 ;
        RECT 72.090 2.195 75.570 4.280 ;
        RECT 76.690 2.195 80.170 4.280 ;
        RECT 81.290 2.195 84.770 4.280 ;
        RECT 85.890 2.195 89.370 4.280 ;
        RECT 90.490 2.195 93.970 4.280 ;
        RECT 95.090 2.195 98.570 4.280 ;
        RECT 99.690 2.195 103.170 4.280 ;
        RECT 104.290 2.195 107.770 4.280 ;
        RECT 108.890 2.195 112.370 4.280 ;
        RECT 113.490 2.195 116.970 4.280 ;
        RECT 118.090 2.195 121.570 4.280 ;
        RECT 122.690 2.195 126.170 4.280 ;
        RECT 127.290 2.195 130.770 4.280 ;
        RECT 131.890 2.195 135.370 4.280 ;
        RECT 136.490 2.195 139.970 4.280 ;
        RECT 141.090 2.195 144.570 4.280 ;
        RECT 145.690 2.195 149.170 4.280 ;
        RECT 150.290 2.195 154.230 4.280 ;
        RECT 155.350 2.195 158.830 4.280 ;
        RECT 159.950 2.195 163.430 4.280 ;
        RECT 164.550 2.195 168.030 4.280 ;
        RECT 169.150 2.195 172.630 4.280 ;
        RECT 173.750 2.195 177.230 4.280 ;
        RECT 178.350 2.195 181.830 4.280 ;
        RECT 182.950 2.195 186.430 4.280 ;
        RECT 187.550 2.195 191.030 4.280 ;
        RECT 192.150 2.195 195.630 4.280 ;
        RECT 196.750 2.195 200.230 4.280 ;
        RECT 201.350 2.195 204.830 4.280 ;
        RECT 205.950 2.195 209.430 4.280 ;
        RECT 210.550 2.195 214.030 4.280 ;
        RECT 215.150 2.195 218.630 4.280 ;
        RECT 219.750 2.195 223.230 4.280 ;
        RECT 224.350 2.195 227.830 4.280 ;
        RECT 228.950 2.195 232.430 4.280 ;
        RECT 233.550 2.195 237.030 4.280 ;
        RECT 238.150 2.195 241.630 4.280 ;
        RECT 242.750 2.195 246.230 4.280 ;
        RECT 247.350 2.195 250.830 4.280 ;
        RECT 251.950 2.195 255.430 4.280 ;
        RECT 256.550 2.195 260.030 4.280 ;
        RECT 261.150 2.195 264.630 4.280 ;
        RECT 265.750 2.195 269.230 4.280 ;
        RECT 270.350 2.195 273.830 4.280 ;
        RECT 274.950 2.195 278.430 4.280 ;
        RECT 279.550 2.195 283.030 4.280 ;
        RECT 284.150 2.195 287.630 4.280 ;
        RECT 288.750 2.195 292.230 4.280 ;
        RECT 293.350 2.195 296.830 4.280 ;
        RECT 297.950 2.195 297.980 4.280 ;
      LAYER met3 ;
        RECT 4.400 297.180 295.600 298.345 ;
        RECT 4.400 296.500 296.000 297.180 ;
        RECT 4.000 296.460 296.000 296.500 ;
        RECT 4.000 294.460 295.600 296.460 ;
        RECT 4.000 293.740 296.000 294.460 ;
        RECT 4.400 291.740 295.600 293.740 ;
        RECT 4.000 291.020 296.000 291.740 ;
        RECT 4.000 289.020 295.600 291.020 ;
        RECT 4.000 288.980 296.000 289.020 ;
        RECT 4.400 288.300 296.000 288.980 ;
        RECT 4.400 286.980 295.600 288.300 ;
        RECT 4.000 286.300 295.600 286.980 ;
        RECT 4.000 285.580 296.000 286.300 ;
        RECT 4.000 284.220 295.600 285.580 ;
        RECT 4.400 283.580 295.600 284.220 ;
        RECT 4.400 283.540 296.000 283.580 ;
        RECT 4.400 282.220 295.600 283.540 ;
        RECT 4.000 281.540 295.600 282.220 ;
        RECT 4.000 280.820 296.000 281.540 ;
        RECT 4.000 279.460 295.600 280.820 ;
        RECT 4.400 278.820 295.600 279.460 ;
        RECT 4.400 278.100 296.000 278.820 ;
        RECT 4.400 277.460 295.600 278.100 ;
        RECT 4.000 276.100 295.600 277.460 ;
        RECT 4.000 275.380 296.000 276.100 ;
        RECT 4.000 274.700 295.600 275.380 ;
        RECT 4.400 273.380 295.600 274.700 ;
        RECT 4.400 272.700 296.000 273.380 ;
        RECT 4.000 272.660 296.000 272.700 ;
        RECT 4.000 270.660 295.600 272.660 ;
        RECT 4.000 269.940 296.000 270.660 ;
        RECT 4.400 267.940 295.600 269.940 ;
        RECT 4.000 267.900 296.000 267.940 ;
        RECT 4.000 265.900 295.600 267.900 ;
        RECT 4.000 265.180 296.000 265.900 ;
        RECT 4.400 263.180 295.600 265.180 ;
        RECT 4.000 262.460 296.000 263.180 ;
        RECT 4.000 260.460 295.600 262.460 ;
        RECT 4.000 260.420 296.000 260.460 ;
        RECT 4.400 259.740 296.000 260.420 ;
        RECT 4.400 258.420 295.600 259.740 ;
        RECT 4.000 257.740 295.600 258.420 ;
        RECT 4.000 257.020 296.000 257.740 ;
        RECT 4.000 256.340 295.600 257.020 ;
        RECT 4.400 255.020 295.600 256.340 ;
        RECT 4.400 254.340 296.000 255.020 ;
        RECT 4.000 254.300 296.000 254.340 ;
        RECT 4.000 252.300 295.600 254.300 ;
        RECT 4.000 252.260 296.000 252.300 ;
        RECT 4.000 251.580 295.600 252.260 ;
        RECT 4.400 250.260 295.600 251.580 ;
        RECT 4.400 249.580 296.000 250.260 ;
        RECT 4.000 249.540 296.000 249.580 ;
        RECT 4.000 247.540 295.600 249.540 ;
        RECT 4.000 246.820 296.000 247.540 ;
        RECT 4.400 244.820 295.600 246.820 ;
        RECT 4.000 244.100 296.000 244.820 ;
        RECT 4.000 242.100 295.600 244.100 ;
        RECT 4.000 242.060 296.000 242.100 ;
        RECT 4.400 241.380 296.000 242.060 ;
        RECT 4.400 240.060 295.600 241.380 ;
        RECT 4.000 239.380 295.600 240.060 ;
        RECT 4.000 238.660 296.000 239.380 ;
        RECT 4.000 237.300 295.600 238.660 ;
        RECT 4.400 236.660 295.600 237.300 ;
        RECT 4.400 236.620 296.000 236.660 ;
        RECT 4.400 235.300 295.600 236.620 ;
        RECT 4.000 234.620 295.600 235.300 ;
        RECT 4.000 233.900 296.000 234.620 ;
        RECT 4.000 232.540 295.600 233.900 ;
        RECT 4.400 231.900 295.600 232.540 ;
        RECT 4.400 231.180 296.000 231.900 ;
        RECT 4.400 230.540 295.600 231.180 ;
        RECT 4.000 229.180 295.600 230.540 ;
        RECT 4.000 228.460 296.000 229.180 ;
        RECT 4.000 227.780 295.600 228.460 ;
        RECT 4.400 226.460 295.600 227.780 ;
        RECT 4.400 225.780 296.000 226.460 ;
        RECT 4.000 225.740 296.000 225.780 ;
        RECT 4.000 223.740 295.600 225.740 ;
        RECT 4.000 223.020 296.000 223.740 ;
        RECT 4.400 221.020 295.600 223.020 ;
        RECT 4.000 220.980 296.000 221.020 ;
        RECT 4.000 218.980 295.600 220.980 ;
        RECT 4.000 218.260 296.000 218.980 ;
        RECT 4.400 216.260 295.600 218.260 ;
        RECT 4.000 215.540 296.000 216.260 ;
        RECT 4.000 214.180 295.600 215.540 ;
        RECT 4.400 213.540 295.600 214.180 ;
        RECT 4.400 212.820 296.000 213.540 ;
        RECT 4.400 212.180 295.600 212.820 ;
        RECT 4.000 210.820 295.600 212.180 ;
        RECT 4.000 210.100 296.000 210.820 ;
        RECT 4.000 209.420 295.600 210.100 ;
        RECT 4.400 208.100 295.600 209.420 ;
        RECT 4.400 207.420 296.000 208.100 ;
        RECT 4.000 207.380 296.000 207.420 ;
        RECT 4.000 205.380 295.600 207.380 ;
        RECT 4.000 205.340 296.000 205.380 ;
        RECT 4.000 204.660 295.600 205.340 ;
        RECT 4.400 203.340 295.600 204.660 ;
        RECT 4.400 202.660 296.000 203.340 ;
        RECT 4.000 202.620 296.000 202.660 ;
        RECT 4.000 200.620 295.600 202.620 ;
        RECT 4.000 199.900 296.000 200.620 ;
        RECT 4.400 197.900 295.600 199.900 ;
        RECT 4.000 197.180 296.000 197.900 ;
        RECT 4.000 195.180 295.600 197.180 ;
        RECT 4.000 195.140 296.000 195.180 ;
        RECT 4.400 194.460 296.000 195.140 ;
        RECT 4.400 193.140 295.600 194.460 ;
        RECT 4.000 192.460 295.600 193.140 ;
        RECT 4.000 191.740 296.000 192.460 ;
        RECT 4.000 190.380 295.600 191.740 ;
        RECT 4.400 189.740 295.600 190.380 ;
        RECT 4.400 189.700 296.000 189.740 ;
        RECT 4.400 188.380 295.600 189.700 ;
        RECT 4.000 187.700 295.600 188.380 ;
        RECT 4.000 186.980 296.000 187.700 ;
        RECT 4.000 185.620 295.600 186.980 ;
        RECT 4.400 184.980 295.600 185.620 ;
        RECT 4.400 184.260 296.000 184.980 ;
        RECT 4.400 183.620 295.600 184.260 ;
        RECT 4.000 182.260 295.600 183.620 ;
        RECT 4.000 181.540 296.000 182.260 ;
        RECT 4.000 180.860 295.600 181.540 ;
        RECT 4.400 179.540 295.600 180.860 ;
        RECT 4.400 178.860 296.000 179.540 ;
        RECT 4.000 178.820 296.000 178.860 ;
        RECT 4.000 176.820 295.600 178.820 ;
        RECT 4.000 176.100 296.000 176.820 ;
        RECT 4.400 174.100 295.600 176.100 ;
        RECT 4.000 174.060 296.000 174.100 ;
        RECT 4.000 172.060 295.600 174.060 ;
        RECT 4.000 172.020 296.000 172.060 ;
        RECT 4.400 171.340 296.000 172.020 ;
        RECT 4.400 170.020 295.600 171.340 ;
        RECT 4.000 169.340 295.600 170.020 ;
        RECT 4.000 168.620 296.000 169.340 ;
        RECT 4.000 167.260 295.600 168.620 ;
        RECT 4.400 166.620 295.600 167.260 ;
        RECT 4.400 165.900 296.000 166.620 ;
        RECT 4.400 165.260 295.600 165.900 ;
        RECT 4.000 163.900 295.600 165.260 ;
        RECT 4.000 163.180 296.000 163.900 ;
        RECT 4.000 162.500 295.600 163.180 ;
        RECT 4.400 161.180 295.600 162.500 ;
        RECT 4.400 160.500 296.000 161.180 ;
        RECT 4.000 160.460 296.000 160.500 ;
        RECT 4.000 158.460 295.600 160.460 ;
        RECT 4.000 158.420 296.000 158.460 ;
        RECT 4.000 157.740 295.600 158.420 ;
        RECT 4.400 156.420 295.600 157.740 ;
        RECT 4.400 155.740 296.000 156.420 ;
        RECT 4.000 155.700 296.000 155.740 ;
        RECT 4.000 153.700 295.600 155.700 ;
        RECT 4.000 152.980 296.000 153.700 ;
        RECT 4.400 150.980 295.600 152.980 ;
        RECT 4.000 150.260 296.000 150.980 ;
        RECT 4.000 148.260 295.600 150.260 ;
        RECT 4.000 148.220 296.000 148.260 ;
        RECT 4.400 147.540 296.000 148.220 ;
        RECT 4.400 146.220 295.600 147.540 ;
        RECT 4.000 145.540 295.600 146.220 ;
        RECT 4.000 144.820 296.000 145.540 ;
        RECT 4.000 143.460 295.600 144.820 ;
        RECT 4.400 142.820 295.600 143.460 ;
        RECT 4.400 142.780 296.000 142.820 ;
        RECT 4.400 141.460 295.600 142.780 ;
        RECT 4.000 140.780 295.600 141.460 ;
        RECT 4.000 140.060 296.000 140.780 ;
        RECT 4.000 138.700 295.600 140.060 ;
        RECT 4.400 138.060 295.600 138.700 ;
        RECT 4.400 137.340 296.000 138.060 ;
        RECT 4.400 136.700 295.600 137.340 ;
        RECT 4.000 135.340 295.600 136.700 ;
        RECT 4.000 134.620 296.000 135.340 ;
        RECT 4.000 133.940 295.600 134.620 ;
        RECT 4.400 132.620 295.600 133.940 ;
        RECT 4.400 131.940 296.000 132.620 ;
        RECT 4.000 131.900 296.000 131.940 ;
        RECT 4.000 129.900 295.600 131.900 ;
        RECT 4.000 129.860 296.000 129.900 ;
        RECT 4.400 129.180 296.000 129.860 ;
        RECT 4.400 127.860 295.600 129.180 ;
        RECT 4.000 127.180 295.600 127.860 ;
        RECT 4.000 127.140 296.000 127.180 ;
        RECT 4.000 125.140 295.600 127.140 ;
        RECT 4.000 125.100 296.000 125.140 ;
        RECT 4.400 124.420 296.000 125.100 ;
        RECT 4.400 123.100 295.600 124.420 ;
        RECT 4.000 122.420 295.600 123.100 ;
        RECT 4.000 121.700 296.000 122.420 ;
        RECT 4.000 120.340 295.600 121.700 ;
        RECT 4.400 119.700 295.600 120.340 ;
        RECT 4.400 118.980 296.000 119.700 ;
        RECT 4.400 118.340 295.600 118.980 ;
        RECT 4.000 116.980 295.600 118.340 ;
        RECT 4.000 116.260 296.000 116.980 ;
        RECT 4.000 115.580 295.600 116.260 ;
        RECT 4.400 114.260 295.600 115.580 ;
        RECT 4.400 113.580 296.000 114.260 ;
        RECT 4.000 113.540 296.000 113.580 ;
        RECT 4.000 111.540 295.600 113.540 ;
        RECT 4.000 111.500 296.000 111.540 ;
        RECT 4.000 110.820 295.600 111.500 ;
        RECT 4.400 109.500 295.600 110.820 ;
        RECT 4.400 108.820 296.000 109.500 ;
        RECT 4.000 108.780 296.000 108.820 ;
        RECT 4.000 106.780 295.600 108.780 ;
        RECT 4.000 106.060 296.000 106.780 ;
        RECT 4.400 104.060 295.600 106.060 ;
        RECT 4.000 103.340 296.000 104.060 ;
        RECT 4.000 101.340 295.600 103.340 ;
        RECT 4.000 101.300 296.000 101.340 ;
        RECT 4.400 100.620 296.000 101.300 ;
        RECT 4.400 99.300 295.600 100.620 ;
        RECT 4.000 98.620 295.600 99.300 ;
        RECT 4.000 97.900 296.000 98.620 ;
        RECT 4.000 96.540 295.600 97.900 ;
        RECT 4.400 95.900 295.600 96.540 ;
        RECT 4.400 95.860 296.000 95.900 ;
        RECT 4.400 94.540 295.600 95.860 ;
        RECT 4.000 93.860 295.600 94.540 ;
        RECT 4.000 93.140 296.000 93.860 ;
        RECT 4.000 91.780 295.600 93.140 ;
        RECT 4.400 91.140 295.600 91.780 ;
        RECT 4.400 90.420 296.000 91.140 ;
        RECT 4.400 89.780 295.600 90.420 ;
        RECT 4.000 88.420 295.600 89.780 ;
        RECT 4.000 87.700 296.000 88.420 ;
        RECT 4.400 85.700 295.600 87.700 ;
        RECT 4.000 84.980 296.000 85.700 ;
        RECT 4.000 82.980 295.600 84.980 ;
        RECT 4.000 82.940 296.000 82.980 ;
        RECT 4.400 82.260 296.000 82.940 ;
        RECT 4.400 80.940 295.600 82.260 ;
        RECT 4.000 80.260 295.600 80.940 ;
        RECT 4.000 80.220 296.000 80.260 ;
        RECT 4.000 78.220 295.600 80.220 ;
        RECT 4.000 78.180 296.000 78.220 ;
        RECT 4.400 77.500 296.000 78.180 ;
        RECT 4.400 76.180 295.600 77.500 ;
        RECT 4.000 75.500 295.600 76.180 ;
        RECT 4.000 74.780 296.000 75.500 ;
        RECT 4.000 73.420 295.600 74.780 ;
        RECT 4.400 72.780 295.600 73.420 ;
        RECT 4.400 72.060 296.000 72.780 ;
        RECT 4.400 71.420 295.600 72.060 ;
        RECT 4.000 70.060 295.600 71.420 ;
        RECT 4.000 69.340 296.000 70.060 ;
        RECT 4.000 68.660 295.600 69.340 ;
        RECT 4.400 67.340 295.600 68.660 ;
        RECT 4.400 66.660 296.000 67.340 ;
        RECT 4.000 66.620 296.000 66.660 ;
        RECT 4.000 64.620 295.600 66.620 ;
        RECT 4.000 64.580 296.000 64.620 ;
        RECT 4.000 63.900 295.600 64.580 ;
        RECT 4.400 62.580 295.600 63.900 ;
        RECT 4.400 61.900 296.000 62.580 ;
        RECT 4.000 61.860 296.000 61.900 ;
        RECT 4.000 59.860 295.600 61.860 ;
        RECT 4.000 59.140 296.000 59.860 ;
        RECT 4.400 57.140 295.600 59.140 ;
        RECT 4.000 56.420 296.000 57.140 ;
        RECT 4.000 54.420 295.600 56.420 ;
        RECT 4.000 54.380 296.000 54.420 ;
        RECT 4.400 53.700 296.000 54.380 ;
        RECT 4.400 52.380 295.600 53.700 ;
        RECT 4.000 51.700 295.600 52.380 ;
        RECT 4.000 50.980 296.000 51.700 ;
        RECT 4.000 49.620 295.600 50.980 ;
        RECT 4.400 48.980 295.600 49.620 ;
        RECT 4.400 48.940 296.000 48.980 ;
        RECT 4.400 47.620 295.600 48.940 ;
        RECT 4.000 46.940 295.600 47.620 ;
        RECT 4.000 46.220 296.000 46.940 ;
        RECT 4.000 45.540 295.600 46.220 ;
        RECT 4.400 44.220 295.600 45.540 ;
        RECT 4.400 43.540 296.000 44.220 ;
        RECT 4.000 43.500 296.000 43.540 ;
        RECT 4.000 41.500 295.600 43.500 ;
        RECT 4.000 40.780 296.000 41.500 ;
        RECT 4.400 38.780 295.600 40.780 ;
        RECT 4.000 38.060 296.000 38.780 ;
        RECT 4.000 36.060 295.600 38.060 ;
        RECT 4.000 36.020 296.000 36.060 ;
        RECT 4.400 35.340 296.000 36.020 ;
        RECT 4.400 34.020 295.600 35.340 ;
        RECT 4.000 33.340 295.600 34.020 ;
        RECT 4.000 33.300 296.000 33.340 ;
        RECT 4.000 31.300 295.600 33.300 ;
        RECT 4.000 31.260 296.000 31.300 ;
        RECT 4.400 30.580 296.000 31.260 ;
        RECT 4.400 29.260 295.600 30.580 ;
        RECT 4.000 28.580 295.600 29.260 ;
        RECT 4.000 27.860 296.000 28.580 ;
        RECT 4.000 26.500 295.600 27.860 ;
        RECT 4.400 25.860 295.600 26.500 ;
        RECT 4.400 25.140 296.000 25.860 ;
        RECT 4.400 24.500 295.600 25.140 ;
        RECT 4.000 23.140 295.600 24.500 ;
        RECT 4.000 22.420 296.000 23.140 ;
        RECT 4.000 21.740 295.600 22.420 ;
        RECT 4.400 20.420 295.600 21.740 ;
        RECT 4.400 19.740 296.000 20.420 ;
        RECT 4.000 19.700 296.000 19.740 ;
        RECT 4.000 17.700 295.600 19.700 ;
        RECT 4.000 17.660 296.000 17.700 ;
        RECT 4.000 16.980 295.600 17.660 ;
        RECT 4.400 15.660 295.600 16.980 ;
        RECT 4.400 14.980 296.000 15.660 ;
        RECT 4.000 14.940 296.000 14.980 ;
        RECT 4.000 12.940 295.600 14.940 ;
        RECT 4.000 12.220 296.000 12.940 ;
        RECT 4.400 10.220 295.600 12.220 ;
        RECT 4.000 9.500 296.000 10.220 ;
        RECT 4.000 7.500 295.600 9.500 ;
        RECT 4.000 7.460 296.000 7.500 ;
        RECT 4.400 6.780 296.000 7.460 ;
        RECT 4.400 5.460 295.600 6.780 ;
        RECT 4.000 4.780 295.600 5.460 ;
        RECT 4.000 4.060 296.000 4.780 ;
        RECT 4.000 3.380 295.600 4.060 ;
        RECT 4.400 2.215 295.600 3.380 ;
      LAYER met4 ;
        RECT 100.575 204.175 102.745 235.785 ;
  END
END wrapped_quad_pwm_fet_drivers
END LIBRARY

