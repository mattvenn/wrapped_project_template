VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_qarma
  CLASS BLOCK ;
  FOREIGN wrapped_qarma ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 400.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 396.000 33.490 400.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 1.400 400.000 2.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 106.120 400.000 106.720 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 117.000 400.000 117.600 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 127.200 400.000 127.800 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 138.080 400.000 138.680 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 148.280 400.000 148.880 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 159.160 400.000 159.760 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 169.360 400.000 169.960 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 180.240 400.000 180.840 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 190.440 400.000 191.040 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 201.320 400.000 201.920 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 11.600 400.000 12.200 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 211.520 400.000 212.120 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 221.720 400.000 222.320 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 232.600 400.000 233.200 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 242.800 400.000 243.400 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 253.680 400.000 254.280 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 263.880 400.000 264.480 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 274.760 400.000 275.360 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 284.960 400.000 285.560 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 295.840 400.000 296.440 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 306.040 400.000 306.640 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 21.800 400.000 22.400 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 316.920 400.000 317.520 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 327.120 400.000 327.720 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 338.000 400.000 338.600 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 348.200 400.000 348.800 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 359.080 400.000 359.680 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 369.280 400.000 369.880 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 380.160 400.000 380.760 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 390.360 400.000 390.960 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 32.680 400.000 33.280 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 42.880 400.000 43.480 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 53.760 400.000 54.360 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 63.960 400.000 64.560 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 74.840 400.000 75.440 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 85.040 400.000 85.640 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 95.920 400.000 96.520 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 8.200 400.000 8.800 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 113.600 400.000 114.200 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 123.800 400.000 124.400 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 134.680 400.000 135.280 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 144.880 400.000 145.480 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 155.080 400.000 155.680 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 165.960 400.000 166.560 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 176.160 400.000 176.760 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 187.040 400.000 187.640 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 197.240 400.000 197.840 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 208.120 400.000 208.720 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 18.400 400.000 19.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 218.320 400.000 218.920 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 229.200 400.000 229.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 239.400 400.000 240.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 250.280 400.000 250.880 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 260.480 400.000 261.080 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 271.360 400.000 271.960 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 281.560 400.000 282.160 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 292.440 400.000 293.040 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 302.640 400.000 303.240 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 313.520 400.000 314.120 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 29.280 400.000 29.880 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 323.720 400.000 324.320 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 334.600 400.000 335.200 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 344.800 400.000 345.400 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 355.000 400.000 355.600 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 365.880 400.000 366.480 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 376.080 400.000 376.680 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 386.960 400.000 387.560 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 397.160 400.000 397.760 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 39.480 400.000 40.080 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 50.360 400.000 50.960 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 60.560 400.000 61.160 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 71.440 400.000 72.040 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 81.640 400.000 82.240 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 92.520 400.000 93.120 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 102.720 400.000 103.320 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 4.800 400.000 5.400 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 109.520 400.000 110.120 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 120.400 400.000 121.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 130.600 400.000 131.200 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 141.480 400.000 142.080 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 151.680 400.000 152.280 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 162.560 400.000 163.160 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 172.760 400.000 173.360 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 183.640 400.000 184.240 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 193.840 400.000 194.440 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 204.720 400.000 205.320 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 15.000 400.000 15.600 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 214.920 400.000 215.520 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 225.800 400.000 226.400 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 236.000 400.000 236.600 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 246.880 400.000 247.480 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 257.080 400.000 257.680 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 267.960 400.000 268.560 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 278.160 400.000 278.760 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 288.360 400.000 288.960 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 299.240 400.000 299.840 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 309.440 400.000 310.040 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 25.880 400.000 26.480 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 320.320 400.000 320.920 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 330.520 400.000 331.120 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 341.400 400.000 342.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 351.600 400.000 352.200 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 362.480 400.000 363.080 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 372.680 400.000 373.280 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 383.560 400.000 384.160 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 393.760 400.000 394.360 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 36.080 400.000 36.680 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 46.960 400.000 47.560 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 57.160 400.000 57.760 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 68.040 400.000 68.640 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 78.240 400.000 78.840 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 88.440 400.000 89.040 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 99.320 400.000 99.920 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 0.000 396.890 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 396.000 397.350 400.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 0.000 286.030 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 0.000 323.290 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 0.000 366.070 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 0.000 372.510 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.190 0.000 384.470 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 0.000 390.910 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.480 4.000 261.080 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.520 4.000 280.120 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.760 4.000 292.360 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.000 4.000 304.600 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.200 4.000 365.800 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.520 4.000 212.120 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.680 4.000 390.280 ;
    END
  END la_oenb[31]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 396.000 39.010 400.000 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 396.000 2.670 400.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 396.000 7.730 400.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 396.000 28.430 400.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 396.000 64.770 400.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 396.000 116.750 400.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 396.000 121.810 400.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 396.000 127.330 400.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 396.000 132.390 400.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 396.000 137.450 400.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 396.000 142.970 400.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 396.000 148.030 400.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 396.000 153.090 400.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 396.000 158.150 400.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 396.000 163.670 400.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 396.000 69.830 400.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 396.000 168.730 400.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 396.000 173.790 400.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 396.000 179.310 400.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 396.000 184.370 400.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 396.000 189.430 400.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 396.000 194.950 400.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 396.000 200.010 400.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 396.000 205.070 400.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 396.000 210.130 400.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 396.000 215.650 400.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 396.000 75.350 400.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 396.000 220.710 400.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 396.000 225.770 400.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 396.000 80.410 400.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 396.000 85.470 400.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 396.000 90.990 400.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 396.000 96.050 400.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 396.000 101.110 400.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 396.000 106.170 400.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 396.000 111.690 400.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 396.000 17.850 400.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 396.000 231.290 400.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 396.000 283.270 400.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 396.000 288.330 400.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 396.000 293.390 400.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 396.000 298.910 400.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 396.000 303.970 400.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 396.000 309.030 400.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 396.000 314.090 400.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 396.000 319.610 400.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 396.000 324.670 400.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 396.000 329.730 400.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 396.000 236.350 400.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 396.000 335.250 400.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 396.000 340.310 400.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 396.000 345.370 400.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 396.000 350.890 400.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 396.000 355.950 400.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 396.000 361.010 400.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 396.000 366.070 400.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 396.000 371.590 400.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 396.000 376.650 400.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 396.000 381.710 400.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 396.000 241.410 400.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 396.000 387.230 400.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 396.000 392.290 400.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 396.000 246.930 400.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 396.000 251.990 400.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 396.000 257.050 400.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 396.000 262.110 400.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 396.000 267.630 400.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 396.000 272.690 400.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 396.000 277.750 400.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.560 4.000 95.160 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 4.000 138.680 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.320 4.000 150.920 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 396.000 44.070 400.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 396.000 49.130 400.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 396.000 54.190 400.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 396.000 59.710 400.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 396.000 12.790 400.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 396.000 23.370 400.000 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 389.200 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 389.200 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 389.200 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 389.200 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 388.960 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 388.960 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 388.960 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 388.960 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 388.960 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 388.960 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 388.960 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 388.960 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 388.960 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 388.960 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 388.960 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 388.960 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 388.960 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 388.960 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 388.960 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 394.995 389.045 ;
      LAYER met1 ;
        RECT 2.370 10.640 397.370 391.640 ;
      LAYER met2 ;
        RECT 2.950 395.720 7.170 397.645 ;
        RECT 8.010 395.720 12.230 397.645 ;
        RECT 13.070 395.720 17.290 397.645 ;
        RECT 18.130 395.720 22.810 397.645 ;
        RECT 23.650 395.720 27.870 397.645 ;
        RECT 28.710 395.720 32.930 397.645 ;
        RECT 33.770 395.720 38.450 397.645 ;
        RECT 39.290 395.720 43.510 397.645 ;
        RECT 44.350 395.720 48.570 397.645 ;
        RECT 49.410 395.720 53.630 397.645 ;
        RECT 54.470 395.720 59.150 397.645 ;
        RECT 59.990 395.720 64.210 397.645 ;
        RECT 65.050 395.720 69.270 397.645 ;
        RECT 70.110 395.720 74.790 397.645 ;
        RECT 75.630 395.720 79.850 397.645 ;
        RECT 80.690 395.720 84.910 397.645 ;
        RECT 85.750 395.720 90.430 397.645 ;
        RECT 91.270 395.720 95.490 397.645 ;
        RECT 96.330 395.720 100.550 397.645 ;
        RECT 101.390 395.720 105.610 397.645 ;
        RECT 106.450 395.720 111.130 397.645 ;
        RECT 111.970 395.720 116.190 397.645 ;
        RECT 117.030 395.720 121.250 397.645 ;
        RECT 122.090 395.720 126.770 397.645 ;
        RECT 127.610 395.720 131.830 397.645 ;
        RECT 132.670 395.720 136.890 397.645 ;
        RECT 137.730 395.720 142.410 397.645 ;
        RECT 143.250 395.720 147.470 397.645 ;
        RECT 148.310 395.720 152.530 397.645 ;
        RECT 153.370 395.720 157.590 397.645 ;
        RECT 158.430 395.720 163.110 397.645 ;
        RECT 163.950 395.720 168.170 397.645 ;
        RECT 169.010 395.720 173.230 397.645 ;
        RECT 174.070 395.720 178.750 397.645 ;
        RECT 179.590 395.720 183.810 397.645 ;
        RECT 184.650 395.720 188.870 397.645 ;
        RECT 189.710 395.720 194.390 397.645 ;
        RECT 195.230 395.720 199.450 397.645 ;
        RECT 200.290 395.720 204.510 397.645 ;
        RECT 205.350 395.720 209.570 397.645 ;
        RECT 210.410 395.720 215.090 397.645 ;
        RECT 215.930 395.720 220.150 397.645 ;
        RECT 220.990 395.720 225.210 397.645 ;
        RECT 226.050 395.720 230.730 397.645 ;
        RECT 231.570 395.720 235.790 397.645 ;
        RECT 236.630 395.720 240.850 397.645 ;
        RECT 241.690 395.720 246.370 397.645 ;
        RECT 247.210 395.720 251.430 397.645 ;
        RECT 252.270 395.720 256.490 397.645 ;
        RECT 257.330 395.720 261.550 397.645 ;
        RECT 262.390 395.720 267.070 397.645 ;
        RECT 267.910 395.720 272.130 397.645 ;
        RECT 272.970 395.720 277.190 397.645 ;
        RECT 278.030 395.720 282.710 397.645 ;
        RECT 283.550 395.720 287.770 397.645 ;
        RECT 288.610 395.720 292.830 397.645 ;
        RECT 293.670 395.720 298.350 397.645 ;
        RECT 299.190 395.720 303.410 397.645 ;
        RECT 304.250 395.720 308.470 397.645 ;
        RECT 309.310 395.720 313.530 397.645 ;
        RECT 314.370 395.720 319.050 397.645 ;
        RECT 319.890 395.720 324.110 397.645 ;
        RECT 324.950 395.720 329.170 397.645 ;
        RECT 330.010 395.720 334.690 397.645 ;
        RECT 335.530 395.720 339.750 397.645 ;
        RECT 340.590 395.720 344.810 397.645 ;
        RECT 345.650 395.720 350.330 397.645 ;
        RECT 351.170 395.720 355.390 397.645 ;
        RECT 356.230 395.720 360.450 397.645 ;
        RECT 361.290 395.720 365.510 397.645 ;
        RECT 366.350 395.720 371.030 397.645 ;
        RECT 371.870 395.720 376.090 397.645 ;
        RECT 376.930 395.720 381.150 397.645 ;
        RECT 381.990 395.720 386.670 397.645 ;
        RECT 387.510 395.720 391.730 397.645 ;
        RECT 392.570 395.720 396.790 397.645 ;
        RECT 2.400 4.280 397.340 395.720 ;
        RECT 2.400 1.515 2.570 4.280 ;
        RECT 3.410 1.515 8.550 4.280 ;
        RECT 9.390 1.515 14.530 4.280 ;
        RECT 15.370 1.515 20.970 4.280 ;
        RECT 21.810 1.515 26.950 4.280 ;
        RECT 27.790 1.515 32.930 4.280 ;
        RECT 33.770 1.515 39.370 4.280 ;
        RECT 40.210 1.515 45.350 4.280 ;
        RECT 46.190 1.515 51.790 4.280 ;
        RECT 52.630 1.515 57.770 4.280 ;
        RECT 58.610 1.515 63.750 4.280 ;
        RECT 64.590 1.515 70.190 4.280 ;
        RECT 71.030 1.515 76.170 4.280 ;
        RECT 77.010 1.515 82.610 4.280 ;
        RECT 83.450 1.515 88.590 4.280 ;
        RECT 89.430 1.515 94.570 4.280 ;
        RECT 95.410 1.515 101.010 4.280 ;
        RECT 101.850 1.515 106.990 4.280 ;
        RECT 107.830 1.515 112.970 4.280 ;
        RECT 113.810 1.515 119.410 4.280 ;
        RECT 120.250 1.515 125.390 4.280 ;
        RECT 126.230 1.515 131.830 4.280 ;
        RECT 132.670 1.515 137.810 4.280 ;
        RECT 138.650 1.515 143.790 4.280 ;
        RECT 144.630 1.515 150.230 4.280 ;
        RECT 151.070 1.515 156.210 4.280 ;
        RECT 157.050 1.515 162.650 4.280 ;
        RECT 163.490 1.515 168.630 4.280 ;
        RECT 169.470 1.515 174.610 4.280 ;
        RECT 175.450 1.515 181.050 4.280 ;
        RECT 181.890 1.515 187.030 4.280 ;
        RECT 187.870 1.515 193.010 4.280 ;
        RECT 193.850 1.515 199.450 4.280 ;
        RECT 200.290 1.515 205.430 4.280 ;
        RECT 206.270 1.515 211.870 4.280 ;
        RECT 212.710 1.515 217.850 4.280 ;
        RECT 218.690 1.515 223.830 4.280 ;
        RECT 224.670 1.515 230.270 4.280 ;
        RECT 231.110 1.515 236.250 4.280 ;
        RECT 237.090 1.515 242.690 4.280 ;
        RECT 243.530 1.515 248.670 4.280 ;
        RECT 249.510 1.515 254.650 4.280 ;
        RECT 255.490 1.515 261.090 4.280 ;
        RECT 261.930 1.515 267.070 4.280 ;
        RECT 267.910 1.515 273.050 4.280 ;
        RECT 273.890 1.515 279.490 4.280 ;
        RECT 280.330 1.515 285.470 4.280 ;
        RECT 286.310 1.515 291.910 4.280 ;
        RECT 292.750 1.515 297.890 4.280 ;
        RECT 298.730 1.515 303.870 4.280 ;
        RECT 304.710 1.515 310.310 4.280 ;
        RECT 311.150 1.515 316.290 4.280 ;
        RECT 317.130 1.515 322.730 4.280 ;
        RECT 323.570 1.515 328.710 4.280 ;
        RECT 329.550 1.515 334.690 4.280 ;
        RECT 335.530 1.515 341.130 4.280 ;
        RECT 341.970 1.515 347.110 4.280 ;
        RECT 347.950 1.515 353.090 4.280 ;
        RECT 353.930 1.515 359.530 4.280 ;
        RECT 360.370 1.515 365.510 4.280 ;
        RECT 366.350 1.515 371.950 4.280 ;
        RECT 372.790 1.515 377.930 4.280 ;
        RECT 378.770 1.515 383.910 4.280 ;
        RECT 384.750 1.515 390.350 4.280 ;
        RECT 391.190 1.515 396.330 4.280 ;
        RECT 397.170 1.515 397.340 4.280 ;
      LAYER met3 ;
        RECT 4.000 396.800 395.600 397.625 ;
        RECT 4.400 396.760 395.600 396.800 ;
        RECT 4.400 395.400 396.000 396.760 ;
        RECT 4.000 394.760 396.000 395.400 ;
        RECT 4.000 393.360 395.600 394.760 ;
        RECT 4.000 391.360 396.000 393.360 ;
        RECT 4.000 390.680 395.600 391.360 ;
        RECT 4.400 389.960 395.600 390.680 ;
        RECT 4.400 389.280 396.000 389.960 ;
        RECT 4.000 387.960 396.000 389.280 ;
        RECT 4.000 386.560 395.600 387.960 ;
        RECT 4.000 384.560 396.000 386.560 ;
        RECT 4.400 383.160 395.600 384.560 ;
        RECT 4.000 381.160 396.000 383.160 ;
        RECT 4.000 379.760 395.600 381.160 ;
        RECT 4.000 378.440 396.000 379.760 ;
        RECT 4.400 377.080 396.000 378.440 ;
        RECT 4.400 377.040 395.600 377.080 ;
        RECT 4.000 375.680 395.600 377.040 ;
        RECT 4.000 373.680 396.000 375.680 ;
        RECT 4.000 372.320 395.600 373.680 ;
        RECT 4.400 372.280 395.600 372.320 ;
        RECT 4.400 370.920 396.000 372.280 ;
        RECT 4.000 370.280 396.000 370.920 ;
        RECT 4.000 368.880 395.600 370.280 ;
        RECT 4.000 366.880 396.000 368.880 ;
        RECT 4.000 366.200 395.600 366.880 ;
        RECT 4.400 365.480 395.600 366.200 ;
        RECT 4.400 364.800 396.000 365.480 ;
        RECT 4.000 363.480 396.000 364.800 ;
        RECT 4.000 362.080 395.600 363.480 ;
        RECT 4.000 360.080 396.000 362.080 ;
        RECT 4.400 358.680 395.600 360.080 ;
        RECT 4.000 356.000 396.000 358.680 ;
        RECT 4.000 354.600 395.600 356.000 ;
        RECT 4.000 353.960 396.000 354.600 ;
        RECT 4.400 352.600 396.000 353.960 ;
        RECT 4.400 352.560 395.600 352.600 ;
        RECT 4.000 351.200 395.600 352.560 ;
        RECT 4.000 349.200 396.000 351.200 ;
        RECT 4.000 347.840 395.600 349.200 ;
        RECT 4.400 347.800 395.600 347.840 ;
        RECT 4.400 346.440 396.000 347.800 ;
        RECT 4.000 345.800 396.000 346.440 ;
        RECT 4.000 344.400 395.600 345.800 ;
        RECT 4.000 342.400 396.000 344.400 ;
        RECT 4.000 341.720 395.600 342.400 ;
        RECT 4.400 341.000 395.600 341.720 ;
        RECT 4.400 340.320 396.000 341.000 ;
        RECT 4.000 339.000 396.000 340.320 ;
        RECT 4.000 337.600 395.600 339.000 ;
        RECT 4.000 335.600 396.000 337.600 ;
        RECT 4.400 334.200 395.600 335.600 ;
        RECT 4.000 331.520 396.000 334.200 ;
        RECT 4.000 330.120 395.600 331.520 ;
        RECT 4.000 329.480 396.000 330.120 ;
        RECT 4.400 328.120 396.000 329.480 ;
        RECT 4.400 328.080 395.600 328.120 ;
        RECT 4.000 326.720 395.600 328.080 ;
        RECT 4.000 324.720 396.000 326.720 ;
        RECT 4.000 323.360 395.600 324.720 ;
        RECT 4.400 323.320 395.600 323.360 ;
        RECT 4.400 321.960 396.000 323.320 ;
        RECT 4.000 321.320 396.000 321.960 ;
        RECT 4.000 319.920 395.600 321.320 ;
        RECT 4.000 317.920 396.000 319.920 ;
        RECT 4.000 317.240 395.600 317.920 ;
        RECT 4.400 316.520 395.600 317.240 ;
        RECT 4.400 315.840 396.000 316.520 ;
        RECT 4.000 314.520 396.000 315.840 ;
        RECT 4.000 313.120 395.600 314.520 ;
        RECT 4.000 311.120 396.000 313.120 ;
        RECT 4.400 310.440 396.000 311.120 ;
        RECT 4.400 309.720 395.600 310.440 ;
        RECT 4.000 309.040 395.600 309.720 ;
        RECT 4.000 307.040 396.000 309.040 ;
        RECT 4.000 305.640 395.600 307.040 ;
        RECT 4.000 305.000 396.000 305.640 ;
        RECT 4.400 303.640 396.000 305.000 ;
        RECT 4.400 303.600 395.600 303.640 ;
        RECT 4.000 302.240 395.600 303.600 ;
        RECT 4.000 300.240 396.000 302.240 ;
        RECT 4.000 298.880 395.600 300.240 ;
        RECT 4.400 298.840 395.600 298.880 ;
        RECT 4.400 297.480 396.000 298.840 ;
        RECT 4.000 296.840 396.000 297.480 ;
        RECT 4.000 295.440 395.600 296.840 ;
        RECT 4.000 293.440 396.000 295.440 ;
        RECT 4.000 292.760 395.600 293.440 ;
        RECT 4.400 292.040 395.600 292.760 ;
        RECT 4.400 291.360 396.000 292.040 ;
        RECT 4.000 289.360 396.000 291.360 ;
        RECT 4.000 287.960 395.600 289.360 ;
        RECT 4.000 286.640 396.000 287.960 ;
        RECT 4.400 285.960 396.000 286.640 ;
        RECT 4.400 285.240 395.600 285.960 ;
        RECT 4.000 284.560 395.600 285.240 ;
        RECT 4.000 282.560 396.000 284.560 ;
        RECT 4.000 281.160 395.600 282.560 ;
        RECT 4.000 280.520 396.000 281.160 ;
        RECT 4.400 279.160 396.000 280.520 ;
        RECT 4.400 279.120 395.600 279.160 ;
        RECT 4.000 277.760 395.600 279.120 ;
        RECT 4.000 275.760 396.000 277.760 ;
        RECT 4.000 274.400 395.600 275.760 ;
        RECT 4.400 274.360 395.600 274.400 ;
        RECT 4.400 273.000 396.000 274.360 ;
        RECT 4.000 272.360 396.000 273.000 ;
        RECT 4.000 270.960 395.600 272.360 ;
        RECT 4.000 268.960 396.000 270.960 ;
        RECT 4.000 267.600 395.600 268.960 ;
        RECT 4.400 267.560 395.600 267.600 ;
        RECT 4.400 266.200 396.000 267.560 ;
        RECT 4.000 264.880 396.000 266.200 ;
        RECT 4.000 263.480 395.600 264.880 ;
        RECT 4.000 261.480 396.000 263.480 ;
        RECT 4.400 260.080 395.600 261.480 ;
        RECT 4.000 258.080 396.000 260.080 ;
        RECT 4.000 256.680 395.600 258.080 ;
        RECT 4.000 255.360 396.000 256.680 ;
        RECT 4.400 254.680 396.000 255.360 ;
        RECT 4.400 253.960 395.600 254.680 ;
        RECT 4.000 253.280 395.600 253.960 ;
        RECT 4.000 251.280 396.000 253.280 ;
        RECT 4.000 249.880 395.600 251.280 ;
        RECT 4.000 249.240 396.000 249.880 ;
        RECT 4.400 247.880 396.000 249.240 ;
        RECT 4.400 247.840 395.600 247.880 ;
        RECT 4.000 246.480 395.600 247.840 ;
        RECT 4.000 243.800 396.000 246.480 ;
        RECT 4.000 243.120 395.600 243.800 ;
        RECT 4.400 242.400 395.600 243.120 ;
        RECT 4.400 241.720 396.000 242.400 ;
        RECT 4.000 240.400 396.000 241.720 ;
        RECT 4.000 239.000 395.600 240.400 ;
        RECT 4.000 237.000 396.000 239.000 ;
        RECT 4.400 235.600 395.600 237.000 ;
        RECT 4.000 233.600 396.000 235.600 ;
        RECT 4.000 232.200 395.600 233.600 ;
        RECT 4.000 230.880 396.000 232.200 ;
        RECT 4.400 230.200 396.000 230.880 ;
        RECT 4.400 229.480 395.600 230.200 ;
        RECT 4.000 228.800 395.600 229.480 ;
        RECT 4.000 226.800 396.000 228.800 ;
        RECT 4.000 225.400 395.600 226.800 ;
        RECT 4.000 224.760 396.000 225.400 ;
        RECT 4.400 223.360 396.000 224.760 ;
        RECT 4.000 222.720 396.000 223.360 ;
        RECT 4.000 221.320 395.600 222.720 ;
        RECT 4.000 219.320 396.000 221.320 ;
        RECT 4.000 218.640 395.600 219.320 ;
        RECT 4.400 217.920 395.600 218.640 ;
        RECT 4.400 217.240 396.000 217.920 ;
        RECT 4.000 215.920 396.000 217.240 ;
        RECT 4.000 214.520 395.600 215.920 ;
        RECT 4.000 212.520 396.000 214.520 ;
        RECT 4.400 211.120 395.600 212.520 ;
        RECT 4.000 209.120 396.000 211.120 ;
        RECT 4.000 207.720 395.600 209.120 ;
        RECT 4.000 206.400 396.000 207.720 ;
        RECT 4.400 205.720 396.000 206.400 ;
        RECT 4.400 205.000 395.600 205.720 ;
        RECT 4.000 204.320 395.600 205.000 ;
        RECT 4.000 202.320 396.000 204.320 ;
        RECT 4.000 200.920 395.600 202.320 ;
        RECT 4.000 200.280 396.000 200.920 ;
        RECT 4.400 198.880 396.000 200.280 ;
        RECT 4.000 198.240 396.000 198.880 ;
        RECT 4.000 196.840 395.600 198.240 ;
        RECT 4.000 194.840 396.000 196.840 ;
        RECT 4.000 194.160 395.600 194.840 ;
        RECT 4.400 193.440 395.600 194.160 ;
        RECT 4.400 192.760 396.000 193.440 ;
        RECT 4.000 191.440 396.000 192.760 ;
        RECT 4.000 190.040 395.600 191.440 ;
        RECT 4.000 188.040 396.000 190.040 ;
        RECT 4.400 186.640 395.600 188.040 ;
        RECT 4.000 184.640 396.000 186.640 ;
        RECT 4.000 183.240 395.600 184.640 ;
        RECT 4.000 181.920 396.000 183.240 ;
        RECT 4.400 181.240 396.000 181.920 ;
        RECT 4.400 180.520 395.600 181.240 ;
        RECT 4.000 179.840 395.600 180.520 ;
        RECT 4.000 177.160 396.000 179.840 ;
        RECT 4.000 175.800 395.600 177.160 ;
        RECT 4.400 175.760 395.600 175.800 ;
        RECT 4.400 174.400 396.000 175.760 ;
        RECT 4.000 173.760 396.000 174.400 ;
        RECT 4.000 172.360 395.600 173.760 ;
        RECT 4.000 170.360 396.000 172.360 ;
        RECT 4.000 169.680 395.600 170.360 ;
        RECT 4.400 168.960 395.600 169.680 ;
        RECT 4.400 168.280 396.000 168.960 ;
        RECT 4.000 166.960 396.000 168.280 ;
        RECT 4.000 165.560 395.600 166.960 ;
        RECT 4.000 163.560 396.000 165.560 ;
        RECT 4.400 162.160 395.600 163.560 ;
        RECT 4.000 160.160 396.000 162.160 ;
        RECT 4.000 158.760 395.600 160.160 ;
        RECT 4.000 157.440 396.000 158.760 ;
        RECT 4.400 156.080 396.000 157.440 ;
        RECT 4.400 156.040 395.600 156.080 ;
        RECT 4.000 154.680 395.600 156.040 ;
        RECT 4.000 152.680 396.000 154.680 ;
        RECT 4.000 151.320 395.600 152.680 ;
        RECT 4.400 151.280 395.600 151.320 ;
        RECT 4.400 149.920 396.000 151.280 ;
        RECT 4.000 149.280 396.000 149.920 ;
        RECT 4.000 147.880 395.600 149.280 ;
        RECT 4.000 145.880 396.000 147.880 ;
        RECT 4.000 145.200 395.600 145.880 ;
        RECT 4.400 144.480 395.600 145.200 ;
        RECT 4.400 143.800 396.000 144.480 ;
        RECT 4.000 142.480 396.000 143.800 ;
        RECT 4.000 141.080 395.600 142.480 ;
        RECT 4.000 139.080 396.000 141.080 ;
        RECT 4.400 137.680 395.600 139.080 ;
        RECT 4.000 135.680 396.000 137.680 ;
        RECT 4.000 134.280 395.600 135.680 ;
        RECT 4.000 132.280 396.000 134.280 ;
        RECT 4.400 131.600 396.000 132.280 ;
        RECT 4.400 130.880 395.600 131.600 ;
        RECT 4.000 130.200 395.600 130.880 ;
        RECT 4.000 128.200 396.000 130.200 ;
        RECT 4.000 126.800 395.600 128.200 ;
        RECT 4.000 126.160 396.000 126.800 ;
        RECT 4.400 124.800 396.000 126.160 ;
        RECT 4.400 124.760 395.600 124.800 ;
        RECT 4.000 123.400 395.600 124.760 ;
        RECT 4.000 121.400 396.000 123.400 ;
        RECT 4.000 120.040 395.600 121.400 ;
        RECT 4.400 120.000 395.600 120.040 ;
        RECT 4.400 118.640 396.000 120.000 ;
        RECT 4.000 118.000 396.000 118.640 ;
        RECT 4.000 116.600 395.600 118.000 ;
        RECT 4.000 114.600 396.000 116.600 ;
        RECT 4.000 113.920 395.600 114.600 ;
        RECT 4.400 113.200 395.600 113.920 ;
        RECT 4.400 112.520 396.000 113.200 ;
        RECT 4.000 110.520 396.000 112.520 ;
        RECT 4.000 109.120 395.600 110.520 ;
        RECT 4.000 107.800 396.000 109.120 ;
        RECT 4.400 107.120 396.000 107.800 ;
        RECT 4.400 106.400 395.600 107.120 ;
        RECT 4.000 105.720 395.600 106.400 ;
        RECT 4.000 103.720 396.000 105.720 ;
        RECT 4.000 102.320 395.600 103.720 ;
        RECT 4.000 101.680 396.000 102.320 ;
        RECT 4.400 100.320 396.000 101.680 ;
        RECT 4.400 100.280 395.600 100.320 ;
        RECT 4.000 98.920 395.600 100.280 ;
        RECT 4.000 96.920 396.000 98.920 ;
        RECT 4.000 95.560 395.600 96.920 ;
        RECT 4.400 95.520 395.600 95.560 ;
        RECT 4.400 94.160 396.000 95.520 ;
        RECT 4.000 93.520 396.000 94.160 ;
        RECT 4.000 92.120 395.600 93.520 ;
        RECT 4.000 89.440 396.000 92.120 ;
        RECT 4.400 88.040 395.600 89.440 ;
        RECT 4.000 86.040 396.000 88.040 ;
        RECT 4.000 84.640 395.600 86.040 ;
        RECT 4.000 83.320 396.000 84.640 ;
        RECT 4.400 82.640 396.000 83.320 ;
        RECT 4.400 81.920 395.600 82.640 ;
        RECT 4.000 81.240 395.600 81.920 ;
        RECT 4.000 79.240 396.000 81.240 ;
        RECT 4.000 77.840 395.600 79.240 ;
        RECT 4.000 77.200 396.000 77.840 ;
        RECT 4.400 75.840 396.000 77.200 ;
        RECT 4.400 75.800 395.600 75.840 ;
        RECT 4.000 74.440 395.600 75.800 ;
        RECT 4.000 72.440 396.000 74.440 ;
        RECT 4.000 71.080 395.600 72.440 ;
        RECT 4.400 71.040 395.600 71.080 ;
        RECT 4.400 69.680 396.000 71.040 ;
        RECT 4.000 69.040 396.000 69.680 ;
        RECT 4.000 67.640 395.600 69.040 ;
        RECT 4.000 64.960 396.000 67.640 ;
        RECT 4.400 63.560 395.600 64.960 ;
        RECT 4.000 61.560 396.000 63.560 ;
        RECT 4.000 60.160 395.600 61.560 ;
        RECT 4.000 58.840 396.000 60.160 ;
        RECT 4.400 58.160 396.000 58.840 ;
        RECT 4.400 57.440 395.600 58.160 ;
        RECT 4.000 56.760 395.600 57.440 ;
        RECT 4.000 54.760 396.000 56.760 ;
        RECT 4.000 53.360 395.600 54.760 ;
        RECT 4.000 52.720 396.000 53.360 ;
        RECT 4.400 51.360 396.000 52.720 ;
        RECT 4.400 51.320 395.600 51.360 ;
        RECT 4.000 49.960 395.600 51.320 ;
        RECT 4.000 47.960 396.000 49.960 ;
        RECT 4.000 46.600 395.600 47.960 ;
        RECT 4.400 46.560 395.600 46.600 ;
        RECT 4.400 45.200 396.000 46.560 ;
        RECT 4.000 43.880 396.000 45.200 ;
        RECT 4.000 42.480 395.600 43.880 ;
        RECT 4.000 40.480 396.000 42.480 ;
        RECT 4.400 39.080 395.600 40.480 ;
        RECT 4.000 37.080 396.000 39.080 ;
        RECT 4.000 35.680 395.600 37.080 ;
        RECT 4.000 34.360 396.000 35.680 ;
        RECT 4.400 33.680 396.000 34.360 ;
        RECT 4.400 32.960 395.600 33.680 ;
        RECT 4.000 32.280 395.600 32.960 ;
        RECT 4.000 30.280 396.000 32.280 ;
        RECT 4.000 28.880 395.600 30.280 ;
        RECT 4.000 28.240 396.000 28.880 ;
        RECT 4.400 26.880 396.000 28.240 ;
        RECT 4.400 26.840 395.600 26.880 ;
        RECT 4.000 25.480 395.600 26.840 ;
        RECT 4.000 22.800 396.000 25.480 ;
        RECT 4.000 22.120 395.600 22.800 ;
        RECT 4.400 21.400 395.600 22.120 ;
        RECT 4.400 20.720 396.000 21.400 ;
        RECT 4.000 19.400 396.000 20.720 ;
        RECT 4.000 18.000 395.600 19.400 ;
        RECT 4.000 16.000 396.000 18.000 ;
        RECT 4.400 14.600 395.600 16.000 ;
        RECT 4.000 12.600 396.000 14.600 ;
        RECT 4.000 11.200 395.600 12.600 ;
        RECT 4.000 9.880 396.000 11.200 ;
        RECT 4.400 9.200 396.000 9.880 ;
        RECT 4.400 8.480 395.600 9.200 ;
        RECT 4.000 7.800 395.600 8.480 ;
        RECT 4.000 5.800 396.000 7.800 ;
        RECT 4.000 4.400 395.600 5.800 ;
        RECT 4.000 3.760 396.000 4.400 ;
        RECT 4.400 2.400 396.000 3.760 ;
        RECT 4.400 2.360 395.600 2.400 ;
        RECT 4.000 1.535 395.600 2.360 ;
      LAYER met4 ;
        RECT 48.135 96.735 97.440 370.425 ;
        RECT 99.840 96.735 100.740 370.425 ;
        RECT 103.140 96.735 104.040 370.425 ;
        RECT 106.440 96.735 107.340 370.425 ;
        RECT 109.740 96.735 174.240 370.425 ;
        RECT 176.640 96.735 177.540 370.425 ;
        RECT 179.940 96.735 180.840 370.425 ;
        RECT 183.240 96.735 184.140 370.425 ;
        RECT 186.540 96.735 251.040 370.425 ;
        RECT 253.440 96.735 254.340 370.425 ;
        RECT 256.740 96.735 257.640 370.425 ;
        RECT 260.040 96.735 260.940 370.425 ;
        RECT 263.340 96.735 327.225 370.425 ;
  END
END wrapped_qarma
END LIBRARY

